--
--Written by GowinSynthesis
--Product Version "V1.9.9 Beta-4 Education"
--Tue Nov 28 23:35:53 2023

--Source file index table:
--file0 "\/home/cod3r/Data/vhdl/Gowin/IDE/ipcore/DDR3/data/ddr3_1_4code_hs/ddr3_1_4code_hs.v"
--file1 "\/home/cod3r/Data/vhdl/Gowin/IDE/ipcore/DDR3/data/ddr3_1_4code_hs/DDR3_TOP.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
nUzstHBazk1VVexUhY/Vf60d44VWVyAPRBY1vK2YhLWlQ+/KrcTN0atIMM9wVYAvXqbex2FeXzv5
gL5etDaWo92ahAtD5KCoK89DnhNisE7fcsOP6ij200VD7d4VqjAXy6x3UQ6mrx2QVQmgvVDUwcmw
M31//3G4qOhjqUqOXE1G3cLS2GWUmp0ff+FJkU5afiGKRLE21rtzKIFdUqlIUY3Nl4ocMuGGY+Qn
Bo/6HmJ3WrpCsAKfeGFaa3HPllyoZCm2fvY00DD4E4NjX7oxKHMT12XGG0hRjFOqSeKBv7ZDLRyB
JIWCwblrRJGeqUSmdLo6oNJYWRxtK/bh481BSw==

`protect encoding=(enctype="base64", line_length=76, bytes=1102160)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
n+rgrt+9g31QvgQfj3knN5xGnkuJE3mh+Egu712unF1deD2bKxy6AonLPTkk6vjySqTZ2ujWIuay
tGcpUQK6ur6xNt4Ml6Xjp9VlmCSvWCKbLYe1fyMjQ9ISRqteIfDsMSenshB+jg+94/09KjWfJvNi
mLY5MShwwUjZBWFUUE0gOLeobRvfXG3zpjamTnKSsv2URiq77VOv0xPW9XK+zukPnibWaPdw5zUV
zfPfm2YH9ty0uY78lB5hM0y0V7ioJFOx1eyPWCkXRBCBxjGTw5vaPEuExvOtbUFyAVl3JsBuzisI
QRQBbKuOMM4KNcDE1Buoyq4xRZTW7IpBNbGobmKU/Lu0B70UHxUz/Ae69TcpfEuPQ/6KO5Yno+vf
0HAMT86IX8AMCYovIn3uGBlNV7nehMv7hW+lYsofjEpZTAjLWYDWPs/sVecnvehdCdmq5CEfNVnY
Yq358AnxTB/tWq/T6FvZrfldBBO59++5mZTcd/0orNS4bz1GIOtZFTTNXy0AedCxsfhbFAhKYGGg
yiK+wWlR2ffMV7XiuB/d9lNpNJwwr91QH1gaPHIqBQjX650HUX8wgkhzDDEd6xelgHU5Ol+X0ilk
3SfX3nKt/CO3d8D8HRmkWcpUoBvGpIGbx+CC7CJncDxWkTclwBiT7xmnph1+TkSv+ToeBGJ9PsEo
4gE+xReqt6kpxAVKEtJyN3GErbaTM9VayRL/6oUhSV+rJohg8ezebj6srlBtlAVkUvp2ikgaxbTm
EMRPbHb6DlbiJMjPLUe9xFJGL50RZfKxrgE3uQygO1Frz/dLP3HgQQVS0QTGfD1+lOX6m0VRLX1u
tK831p3qu1J6Y3tfwjI5jzOJLMyAvNPZbkHnfcnm4k42OiZbK6oLZO2Q25ExiH6fKHhzNi8Pl0X3
FyWvemoMsM8I1TCNa7REKmijgIlnhE9q/WmAGmwMuoL8vo5zWmq398y9gfd6VyDkcnvYC7ADO81B
GQhaZ+mLZTwjXdOy6eGGqQpX2ksbEu5s8Wkv1TSIYcS7DXDqQig8bWp6MVhkxRcuUa0zFsZKNNPw
+AXb8VFG7/2jDFftMlDVFrEwhppKgA6G9MLbRXUnbUxrsHFKUp+N2yNJEh8tADG+5gfmRctyXxcU
EdbKbQOSy8h2QuMo6WkHVxZlqQEIzvfVT7ozkUClAX6vOLapvEFLOGCxsjcnxEMw3+kM8rDAdz7q
JxAsA2YFYMWwgjLYgJHOsoeVGJJYQLQic2qi7mO1tgbZh7VexkBspHuf3cUR0ecz07wAI7BZE5qM
YUwkSGmtTmdBygJYSIps+BcKnPBd+dZ1OSCglJlySqJBEq8cD4l4XLNXAlFrHdwxdR4M+OpxF/Y3
U4ZcUByDoUTEU4RX9AtA+9VStmCjMM2Lr3wF+ZVxflMYL2Z3kmtSODzYD1rrfoIFed5K8Nz5ITT6
ZlzGJqnKZRQVJkkNsV/1DKJ1q+zRnvzOYWZ+Az1E8vhL4CF1BukJoLK1q8hiLc8+/JcQ1zYNTg4b
c1pk4UdSYXEqXq0sUJ0bl8OXWjJKHeQdcwqgp3lOkjKRj5GYp7STrgxLFPxRPZKnws09kBjTg8Bs
dsupYyo5yRMxJQMpmoJx9XLU7WBjRYepC04xWy8oE5P4W2UVN2SF375RQz4+kRNlx7jys6SkOP+Z
Ze1yKJHPIT4VLa/Q48BFmuEC/h7UBVk5jy5+0wiePY6P4ZT9wgyqs1xf0NpRsLYMQzSXIiGr+KLh
9TRuro0WmsDFthraOLpXMnO0C9guw6Qdk1I4lzoIkDWmWy83lH60eXwspxXK9Py6Zr/vSZ1zXZmN
R11ASdw2IKlbpqusyAlkD0bTpz/hCeUDDuSzd8amBcgdtuSrn9vAoOtqmKb4WiUuI2rNlIheJYJR
jtFLAVlk6kXpxWuiGBs6NUYSh6+qY7xb00rG4g++cBrLpVYNIPiraoi/KQ4+0TTPDdQaz158JbPl
iwgammZL/eRVwl44OYg1fo+hKm4n4pgAiATAk9hdPieVB55uE/TAxUo+tjAkWI0KENVAzCYxZaWb
OzCL9SzopZeO9GnhZpma3vPE34GbuYYJe1Xeeoh6v28/NbpvyumgqBnYGLUOu/oI6Q/HL0tJuhpn
GACsYAdYP2iN6FPXOruVAX9UwsULNRvOHLxG06l1GSH0Mw/Sugj65NBFh7ToFSXY9fKOwe1u7NaT
Ed1JAXmMBT+vbeLW12Mo6bbt/pp9K9QW12WkB59w79qlH2dchSiz7VribtAG5i1jQJCdvZjxskpH
ooYSc48GmbXeK11TulzQffcW3BerX4my/nDsKgeWXu7yKOTX2XH+HkBGruBCz249FHeE/wuNBv3P
zL3qsxKxbBHd7kuZaSwydJTXgWZAZHUEVVzHIVu5+wL142gGrAi/IaNsKL3juBhJG0yAcVelrgxp
PgingNLCiL/fnoePqlca5YzdRebsspz4AWH7qFL7JFAt/3PMERbsHoHmnRslDAeTFbjNGWDqUBA4
7zimEBOR6WiAo+rTddBbd4WEZYQrrpDuAgNmx8tkij3igetx1W8WYbi/wCWpTGjum81bRnhoFgWG
3tJ5VhwZUpmRhdwC0zqAxB0KWyqdsn//FIuRHS5iLDJ5UfwaUEb0JkFbS9gfet6gEStN1XH4pAUE
41j1bXJR6vsAOqpnKYNU+NuRd0ggw2v8hMK2SlQfBt6639s6NxOZHVVNjewsz3h4W9VoKnrlCas7
CiaOwCQW5+a/+LEun8kVjZk0q0MloTKlGC8gmA77JwqeF8Zf3L0gzCuWIDe1VIjB1KyQSZALlM5L
m1xulAAqBoYL6ThG7dYCilatKFPap0f++HEJyAAy5mPOUrTrE9BFKMXA6csqmrb0a1IADKTVYZnX
7uv95GrqtyKguGkrZlqWq0uRP7PSdqrWujjAA8FecnYn3Hop2SEmG42eZ5AC1+GMfQ5gyLMPloXY
JVTwbWUP9rkodC6aMDoR8Q1xIV/M0LiRvUuJsBzbh9ogJd1rqDX1J0nmiduYQDV6ioyX0lp+Lu/I
lhlCGLBX4VclirWtr4nVL19DgoX3AcYJVAbapJnC10L7T06+1giOtpeRzORWyXkZtALapCqs8fjD
chHY7fOeF1bRY1nHDj3MdTqO3Riqv9u5Pol1YFuvmcOtaCmEGjDu7OAzfu6M/eqohyjs4ri6DjEv
/mnpNDGvtPIKmAodZTN7JbUUGdcZLRC84ImuvBACN/2y8r32nRGj6lwJZeWO4ItSYJuDQNlU1oO5
ZtNzsMbpCM3fk5FIxBtQrwRHdiCu8WgtcuWHDcJE18yvV6Jkc9V4UuZnjLSNf4OCBzm+pdDZF3H6
Eh83kj7PTBaonAwjhV2EZ9HniOdQ7hCGcD/w/AjuCVEbsWkYl+rfX76AA8l0dc7pMqAAg+S+l/Dq
C++HZ7hzlF+WmwNihiue5u4sDPdOHfd69epQcKqJ9JmY++4pqSj6lNuuti4vANX5RN//XPwxBX7L
oSyqij89P7Wtk2ZcuKwx9lC8/zWDepdBOqaAKHYpif/Fg4So58st1IUd+ikGyHj0Oi2Mj5uBhCds
H5wNY3wP7W8rB/0egM1cEE8PBPNnHRb5bsuWTxAI7ZHp3w3puDbnWIrXVvoIfbfdIF4dt3K3+ypw
eODu3+4YGGzWPyACPaP0nvuqv4NpnOreQAoqr23YRl0MgGmClFQN1hPJcJLP4Bm6ZP16A8yqClLK
kDxj5xNyzJhvAhjeyXbkBk0ypdissd1CSYBu3hh9hEBktcvEu2k31wPd8L1AUhJ1bzRc+fa1Js7B
dGUuAPE2+3zUnILwEZp13bECkzhj7sIzDuZxFN4KqgRbNEw9PPox8SAEztimOejv00gUgG7VbWM3
kXhfa6z7lkh0ecnTJAk1MTlqeepUFAxSl+P+30E6qqUJmnprBYe7NVNLNzawdBMHmaAc13wyJFEU
gepIBnf5S9oR1eMu3eLr1GGUlN88o5Ep4pj530b5DwJsiGOWPSe/T3+JqY/Rsq+dDVN7SUP5x+Hd
i0kVsaqzxUdT2Hh6MPEBMJC5NUMNmDKiCtXB0ox2PEYCq+JLOgKda2u4Rx1p7mVlIRhMSw2LaiOd
InY3vf5vZ7QlVDQ19/D1yn6ka7hdkjmQAXlkfaPGl5x2j1a2gQgoMh05PAkUD7POfnkG1OrK8gUH
Yjja0eq0sDwXvIOT5TrMWPY/QVQkwxQtjmXGMuB14GqmOvXl2ZqyUXMnLZQV/Rz5xkd0XEfdhnu2
IlKH3ORTfwz9qtTMB4l1NPwK105mDY9Evqd1Zy1YdUsJl5oICetdUwuWODJfgz/SECP3Dgc7v/rS
1/SPDNkm12SqYw2Apv4HrHA56UbfVCKZNnwutp2eqsnjV0/B7GHXxYevZTmceUOsIyIlsF9pTs0v
6OXswW/PuC6ZSvJceqIMhGTnyW5D2c7nVZpKPkBVBnTe7iDiss/o+5WRbmrRwl7/whyzS3HkcVyc
3RvZvuH0cZpsibKrgSW50ExSIEcklmSM3wcL67OmsZhEH6wnEH681wvhLJzLARPMMUi8LKvwq2s8
9qU3MdgeQFr+rUmJxqURV1cXyHZgNOEqfG54hVz1DVM0LTqRAfrxfx/+/PjYZZM2eaZ1G4YxkkTT
G7Ce69i9DhWeKYxonDjRDqQjHoBpuGDOYOFluENbc0ycsqN6WulRuRjaFHhUUuQg2hj2UGMpyIFU
0XDR4jZW2dxWByOXZa/hQFwGJcpVEBDnkWW8OVb/2Q7dPCfoVLjzV4M/dPHpC+5BlPXKKByVAaiV
A/e8l02TKuaow4gZKPz8QWaQk5Ihx3/SzaTdiTUcIPa0S6MnbcxxdsoojpHobHfiZiHNaQ981Mr7
L9lbkQUd0fqR9SqX7lXaycFqv7Uo8/5kWTUSLlVkJwOjbg28MzlPiqRaKhVwkoJ9B3dteVRyWa47
odZKPLRO1p7Xax/6eRvx6X3XwpwVZqBpSxv5g0skd7YgqDGddyQZ7+VshyKjwq14TbSLtk8s0EqJ
M8oGIje4E6PR/Vyn+/WeE7QX3eRu/bDsp4Pz4cPfOERu/MEDUiDreC8IEw8Mf4iBmhbrTJME/x6F
pIs1qdG+8RIwLzZSG6Dll+ZE8CPYgTcZ8Ur6MW2RzKVASwRl7OVsQcsQKpBeEnOTgDSSD2CLclDu
a6KVRex1PHrAh7U0SJteIpVUhwFO+U4wb2RhaP9mJ1U32AYbwFIZUiMV+B6Tzz8LVXZJ+Vr1fvZT
Q9B9KFT+CFHRPYeSfqzCBtRZLjL1AV93IzgrNLi3xNaq+/ng5huUsWLTOg4/gD37zEcNg8OhoGRf
By5rwmMmkUj0gh90vdQdlzyLFDeSsMZcGpI0CVthdAG6/YJQYaVZCo6abHvcaQIcNqgPoZQ7pY9r
jtPtpzMXv250JeU8Gi+M6sVQjAkOQGqW0H4HIHp+v0EREHWWfbbgeHoL4nB4Vydu5POr+68upI1W
Sqb6v+jrrYGOdieHmULZhBWKgoPNQlXo6OWx3Y2ZvLHiaV96rTxtLibHz8LBZY4Pp4zuTIx9+HfO
PFYvoInoKnLP1Qz6A8dfJSq0ALCNGxjV1JOkWOsx255dYlOJQUW/1oJ4X36VSfI0ffgJ5HIOOSxs
kh/ayHjvuqua+Yd/RCBggM4Wxj0k/tPKHYPvdrTq9DP9QtNTZ4fGSx+zX64dFZ9YR94YgtGjp7Kf
Gxzh2yP9gkYLNOpdeUMXwXK1PfFXaZlfQRF6rvVhTmiu/g/RQ7AJeDJeD1WFGSGsCIhfmOcHKsuS
4JbpUqKc+XZ7sXXNClG95eMdi4m29ay1f9Xzwmmx8QWLGsvZhWNWQeZuYsSDXyUdtgGKO0IsquVk
AqgBZ9XHNXKwISyjGJ6nZsTWy9I9CY9Nin4uEzPiKLUuU1DhJcVpXFYTzkvMtahI9CrkGbFzpgRx
06rUf5x1+L70LWrl+PhlTJYwDToUiWdsolN4R9MTrL3CJp7lTCyJF+Wm2l5eEnwhYzvY62aC9iR4
G860TWZ86polKSm3YglHcMXMZ2K6tb3Oxt5moKz5sPbdEBv7i2xWVFf/hK9IpKW2bC4jy7JI68gK
QE1abKFd7w4zjKV8V4jCQtvofQ+Q5QDDnO6vHbpJ49IoQYKeT+T8RgQb3JdzvLoQy1ckV3ZC7twQ
etWJeRBdPloSkqG9MuwOUn58+qbY97lW8+aIhY0OYf4XVsB7fXaO+RB1MxSf4gInJw11IfNlBQM2
Yvd3p76BorER6m6aOMyOdR/MKCx+y3T9RbfJ65/KydSvDALmxIZI8roYPIsbe63B4aPRlutBTBV0
IV83VBD7kELV8I7JAR9PyBhDnM1TUjkX+HMlqFAsnlh+Ru8OvkOWsaVun0Yf4O3HH1wZCJODmFzd
ddszRahE19ipm1jU4++dxc4l6u/L+fD/BNvlsnn0SqqF2UHuZh8/1g0YgkcwTx6cT7a6cm3ohU1T
DvFTUQqXYSktGabkYI3CB2chp4U7M1HN/FUHNeUd3wjIt9hRWlcwysr5HDnvOLeOCuX7vksBT6AC
bQEPYvkoIcYYKRcnp8ExHSb3JyPol91fAe7jf6NSDm233ru/qbB4D1z9oOdNU/yY/yr9dmg5VqPW
hmKhx1zXSyuA8yh0JA9drSyIbTX3WpFcHN67cgYHYgGa8E8+NcAd2Fx76spBD4g/IaB5Si/ztakX
M/E+N0wL1xwII4QYwEX92Geu9H0fMv0+WF62VIGOZdT/dn608hBa1/B/e7KaVEai2xwarqHMI+Jr
PxBhUBsMzN5T1ZH7hDNk6mlYar21k8Oqitogj2EXzzEOs+OdnQma8ebf5Hiu8WopTdhdLpQBBa1h
h2P/t0pSI39wLEmNMWXt67wu2VTN+82HkQ2Iko6KezL4xMEfLPDRj4bxMBIkQLCA4v3QgQ0h76fY
bhGcfMQ5IhT5+ltFB7YBP8rlPZf1XykLdTY9OxlX9YwAMcLB7TS+6H3P5F/uxZZUaRysfchWgsog
GdQ5t2f2GAKHczxeZW9BeCgC9f+gwjzAzZ61r8czBBXEE/fV9p1nFPATQwPBXQsLTOQIxiPkn6/F
wOHl6bTU4z+YDvlq/OVeOJXrUZUCVkCbVNpA16pfSbw9ieVhn6QTFlAOdb0G3qudArKVGmNeG8yf
41Ii8K6VjRilfoSJmV9BF83eJH6GHRyH01jmiEX1MWRMwoyRfju7xl4sUZFZqS+z7uHw6RsTUiqw
TEYDBHkh33kHhCUpIEkSW33KsfKZjyFfMsAvNHAAMRa2GwT2qCCLCk+FqL0A3ykNBPdU/ZjWfaaD
br2c2uMpEtNfcp8ky6ApEmAlkSxy3dCD/jhayOipFtcnqdwP63jnQVenyonISdh7NsQmwGMY2sso
xJLxtt3YyczvZmxYxyVZnVpqdg92DH4M1TXN20qggFz3QL+E4jvyteDeJzlVcjIUoeCOYoKXVWxR
KfWBqI2DUWySm62n9SHt1jcYkDXv5tSeo/mhr/fThYaPve0dPJvMPUx+dj4pHzYFef7zbjp0p6bu
T48JHgBwRLDyWwrHvS7iFjtkH6EXcCH/eRHWqmexVQ/98EmrUP9PlFGxBAug/zSsDKH0HhlNqWbs
p1zol5eAxe7p/1+ij7DWIXiNNui69GAUJpbe2XMGqJnWHCBrIEFigeR3JicqV8EnKzVg2R4iKl+M
wvVl4YfiaeVNmQUx7L1hZct+OA5+vus+EGTfqYCtR4s0PXTaCeuDJXykH7cNoj+y8RyfrDgp6qqo
LtqE3+c6svUnnFtPKqmk++sCqNADfDzZipEeGOFhnuPPmOeAR333vPRgmoQsY2UATOfYyGhWhIsV
5zloB3BiEAVcNwtL8rgQsT0FHTx3m+Nw8MNr1a7oOVM3qGT0GsdDO+WX7mVuDdaEWaU5eME3iNvG
i3E9ywwC9WZdiXheOCh1+qYyzDGCbSDTo6w7Nyp1WRp3Vv/RGVd2R4Dkp/nFJ0Tlgu4LORxzDFnQ
25HOR1VfcR7Hxu0OGwmLnPMGV2MBO09e/EMaJiJNzGJ9Cq83OZSnHEsRyg5We2D93OSZ8GYix0PY
15g8sH1NIB/Hg/VQ4/VoTfhLFMkXmvUV6jOWP2z6SxyzFiRAhgA5JEQ1CRLjVzLY8INNKMnZA7Jz
GOqWHlKOkKVx3kl4664y4F39V55O0XA3gkArT95oi2L46bDMDY03xecne5UEHk7YZXpSMIZa5PF1
HIE/e36trESTS/kjoc8P68LOs8SomH9fIJSt7/iJL2CiWS9WkxZtlgy2VDpxWJddeNcvCo7TSRwJ
zTDRUiKwjGMCCEqXx3rIDAyXePeTtyy0ZzSa3Jw9U7FP+Z8N7rCrF+0InS1/DTtInXm8OWRUMHCb
7/mnufXbVSOyDQW/HNUpoIzzSbITce5fWx+x89xmvMl+vuXJRsrc4aFVgnCEsDpI2oh/bBMz3ljX
bxDeiWD42KBSoqOSBp9rZ46fx38Oe9oTEWT46wfeQhIGr4MlIr8sUt6MDscVQnooBerwkvTj+YgP
FAr3x+QyyqtRuzw7REum4ZtzqnUlwOa6H9mJmLWXGCKhfWiI3+pfHKwb4Z1TieN0Ffg0hFvuMXKo
pfKc/smITgH/8BI5gzVu0tVJZsMofi6ls1N7PQN92E+hrk31R+kj6ceAGTVZ3bXuqvGHk+htFTHe
te9lXOADOQfRAnhwHxQVMe0V0115h3pue1YNtfdugxhle9cN8lMP6UCwE+vwpTBiJzOkYbYr63dm
LkmBN2wbMygkGuIGOsuX6hLD2AFNJ/6YXro9egSS3CdJKjaVAkRECJz8ndSVRJ3eA9BiDehkGEHV
nXJtkdGK6zihvQGlRA0I43XdD1JrAXyyhvyyBmGkbNp7D9tGKqAvqrqhNsPlJ/Myrl/RblxtFqV4
tmzJb7mWDsvN9SAgq99EJvymyuesetVA1bFWv3bvcrxld7MDQ72h3P8GRkwFQF0y4SEnWDgJP9GF
bdlnfuwCT2LR28NKdujkQw3HoFESkP5p5cfjl3iHBz9XgRXv25JvozFdHgw4WwuPH+J31NGhdS0O
0XcCGwh53a8okzKk8TDFaPBFZ1EWefW6M/kHlosFmI9nGsa8ShTPUw/JDJlwUOHz93ZoijLpEpl1
i1+eO0h6qn3hX8tt7du9cBkl7IoD2rGFxR/gaBA6HNDb0kqFDC5pn9c11QPdexCKmM+eRaaeo43t
n+5llgKxK+yheUPuHYVWLwbjE7eydG9/QNSZYw3S+liNwgl/s2pSvgATf7BYHCgCy1rQ91PEl1we
zHplu8wwLT1Kzu/2guN0zPUwglBXut+kjZE09fyZPGKBC8fxiWo7jYEDZlZRiIUQovdKMOqVrYfk
hEveQGgUpAb7mY3GixXwV1e964QdUOWpZN2rF6gu3F66WPRNi4n4LWRqW1Nokp2zuS18FZdZaOLk
utzYwkjEd6f1+IjIpZjiV4n2leiaaEZprELwV+vHBz1e65bJpDuZAp6K+xdnDjLoGrDzGEHdXuJi
C1huYiKP/o/CyfUyhH+nlH9Ud5cxV69TwiqKLFnsHtcQXcu9UjN5zehdb6+5QPuyUXtnnR+luKQ3
c8/ALpFCG3bXIMbg/Va4N9alJhskiAOU+L2Jlgc1YIMcPC4jYwy90uVz+fGenDSomWCg27Wj3KcB
eO3lAN/ieqGFgJNXNJE0ZXEhOTpKTxrbPX2sVXqn8jw08ev/ODsU5F46F2xaQ5GwGwCG91ZoeYx3
0PvhLNZQdHisgbxcDsCd56wf8Pyd6XzJIYlhQ2ktevQ/fzQrkzE94CpWMoTZBff/UEwUq97SeGu6
LN0VonZ0ooaCz16Qip5OaZCQQEsQ0B3zmoiZ63V+lD6FnuHStKnyW/urvA+1UreJnltSBTfrNtH7
p4HcLVLDlIf/PJ6qH3pXN4sjCl9HFIGBA3grFGllZ0dftmA2u9Vx6ZNufuOm0hXojoBnSMrEde29
QlxrCY39Tg6nxhnNs7d/1AATdZY1VbMQmyDgvaV0sDzLo+vbtYBIpcwVv/+R9LJfzr07EZNps+m/
xJ4n7k1Z4lPghJvomgZ6nZz9LmsxmSIjGBljDwwlWNLBo8pi+gzTpRoUZCG/2PumCPwezggVc6fi
vB3W4Xcjy5TobBvFlCq/sNA4qesZw6L9Pm2AxAKC95N57n6FVRy4yS8CmSQxCmVIh7W4m9xRN2fm
sF73qMvTLCSeZ07iUi4IBQzduEYQGcEC0xtRzRHqlsNCv5i4yRN79z9R6QVKxt46Xh12+XjOdrcD
NdL+57dh/XON8hDdETvLe82n9Lqs8B363Cfl/XSUvxHIr8SNVj0Q2YeJxS5DDNQRluskcRBdH5Sm
qOpQdtrKkTBKiQ+3plFt2wluAsTde421SDjZ6LOyrGdN0DLedOCwVo+bw8Jz/GCVlURtV6ZLXH0k
opbHrzpmklybcnk5qki8waFgHerpT4ZcWUWHWYtGcDLxbEIW2Tsnm0WtQjQSPF+zGv7ZLX2BqORd
UrQL8Bet5nMKILv8/Qh913eUcoT2VnERroVCjPelEInjk8Mj16KVRHSeaVCRm1kxnjL3aVFr7koh
wrJRV5BTO0JvVbzNoaBMDai7pKPoUlfEVPvohyheIXKixyNDh+Oofi/HU/1hyCetnJtJgy0HGqY3
Crr8cwk0uiR9eTWi9RoPB2KsOcF43WowBDzwhLjrA/z5dDmazKZ5rupjE2HqCRS4gAY2OcmopS01
WryKuA5yn15eKSSEIzYdWdmG5r8PIg/nd8bWPwPZj2kqUpJN3XGwEXpAfNcO8wP+n1JX4hCm1SVH
0TxE+Ev5LAXflL/y2aRelPG1ALsPFDezD734fW4mTiXXSHqS9unAOW9MFM/9tu96pu6+eMMsNC7d
SXYvJOvhZWCRH571BqTriEvYbQgp5nCDOKNTkT+F5DfJOXfv6Mthz/Kpozm3cI1ftYsnz4b92yfb
JEFK2BHufjVbjnk7OMeZd+1Hy1DNnSlMicwowcJRVmK2TEBCK1OnGNi3JTxN+lb6FHhu3UtuRRAy
z/LSVGFv/1yo5rDK00MeqGTdZBItdCXvytoizP8Iz/vbDAHChpktkSwgJL595tOX1LTltgEszDEP
pup8nAcMGSLR9M7Q0vf+M7MLgHbaROkBWPUmaMKgGi16cHNoBowTU8VXDm2ZnkXeQbUFFD8zTX1w
UR31qXQC+Xb4saa6Ke8uEINZ4P/2rAsAP+9XPiyzvrz9E9BgaEcPRZcY7HY87vCjlYO+TtQBplhd
fJjrJkJNoDvwvklD519wPr54gFkdYVkeXIgr6JV0js880auKrI8c0j/xstsnRjjUjNOr6QK22+l0
U2wdbkc6BShjQKn5cUZXnjZV6RinvbdODAvmzVaaCCdAJCVZFZVjfb9cAZzuaL0ASTAMj164M1MP
TSP5vyrvAP3v1cRxvQxMvK7eotN3mkceuD3Kx1bropt5u4A+A42+EaJQHqim/tPcy6+awmUjPAED
5ru2HZFZKryU6Dbq1U9Avm4BL7L3wrC59edl3cWv/Bk+h3dtqjwDCeCsUSH/nDy8rMzWBLhXL2/r
ExorVDAFcvUyojy1WAe8TpLlN/Fr4+lkD3Us9zM3hlurZwzdo2gcTs4Oi2OtILCHBQ2xBcnNriss
URLXU4lMPUk4JCA7ju3tAHRBC7vtCNuxgJev8LfSDKe9aWUZGg84UvHmTlRy2ATsidakCHFpT7iy
3/zN/lMV+sSh0kQlGmBb3h4JKGgBcdFxFa+cCxNwMDb2560yCPNdN3iJfifXxSoZSZ/ER2u9rM0J
GPp11iDdxuw/SHuhB9hlVfqsiPkZDcmDFVCXbnniCBGk0H9V8nRd8TODL45A1aLmlLvksljHel6B
dyMXwUHA04xTySxBvVNmiNegDVknfXO+hfac0zE9EehphqK6KY5Ke/MWqIbRll1lHg7x59hhkn4j
CF9x7Uf8NWH5XN/CASA4LyyEeufQQIDeCvzsrP7O0/3fqxO/hbE6UXaW3hP9P1d+YibpW51eMq5T
Jxlbex3PncASxWKWO4s8d/rN2m1S54zwkpdvgZronXg4/BlaoFH3fy4ckzmMk1KLN54ek8ccDQeG
g6xUG1D0LplXwfJoVuGaGWYHeSKc7HdevneaAyNIBQRNMtDwH8K57M2txW/hX9bMOYWvHBfNNwvw
f5q7AT57guixbIn+DE0rKN6bUZajl3ZLMg9s2bGtnIt8q6xBv1xRtTyaRxmSRmuAUUE44nGpu+Uk
qAsTOLZwnhZ/cuQ0L6G2huVB7PZBQU5NkOqbB13G0KB0/ragEH/Um0vvtdutJBHq4cGynANlwKnm
nnrSN+Q7KcL5Temrv3gHlHoz3h7f5TeujKGN3cBp/tq/L5/SFhoDcW+ox/8bE//D8j3hp3Itute9
IaC1y34CiJafe6Iy1CAzessFNKYy3wNbHWIjmlvZUocGwZ2mhazWGdFNa6At97sooX8mCA4iDiw9
phpcqVGqeSBQFhXOHGroE9GXRGdergl6Qu/XZwjnDybgraa0af4cxMFIsBM4e+zRNnPyi55PlrDV
mtTXy11MK+VkwKADHcund7mvjsGy2rjMfLtol6nTEpjCaH15X/XWbCX9n/HU1TtUKVgSkYXOIiWG
A6NgoWCwH9veP17nbQjhIgSG5uEHkLbcZVgeLKMKzf87Qa4AiH6/+iqwIAZFFmCb4DWfv72NsvSL
pcbTXKx65EiSdpC6XDac6ZPKnw3ja21jeft3pLnz4fJRvBdJM/Orxhz8sagkIMxkfv0HNXVON/J6
/NAvhWxps36k9nWTZZNgpUD2SvQxBM44m7QXchTqWvI6sKbWBgNO0Natj+M/IJ4VsUdm1Fnpneud
vJKMkIZRy6jeExKv2jzfgSoHsDj2iE1CDkCd0/9LEvNPWEtdzaIAfzM2Gm3qq7F5vh5GYGt9UW8X
Gn9j7D7hWm856UrWx4kM8lPckdclZZyWOgnb4l2fJdK8GG9axQX6A2t74TvDAz1Xay87A7YTAJX+
BHc4d6y5EBpBz2ypsES5r4lEu4m3q/kdkHgHNkBnkJdTol6JV01Sn7RJqkgSF2ZM1uWD2ofX3Kms
LOfm5sCBhuJnSymeQrLBrhxiA6O/M1OFYEJoe8AO5dsPRzVqkiXlkbRbRDao0AtJD1a/f7FnaVlp
qxmJvacRyDLtWy9TltctHXnQVi0lLTTkDziyJUEZjokIpqMAd0v7cfkD9rdpxCpCwZp0ReUyA4j0
TU1hLh1xK+jW9Orhj2tFv+DGvYHX7UVNNJR72751gbuEIGhE3kLTsgT+fY/XUIDR48Iqs7xVwvx0
d68JtwaO8Owtn+YcP0GB4tdq18M+GWSTveLt3/96+x6gokK3+pFPBfQxS6ECKUAMjNPge5WhU6vL
NSgFEc9ERfc48k0TZD6/w6riWd30ZL+wBV/2ynUCkn37qFE+yl8ySbFwTGgmn2O0gE++Ubs/qKfp
qI+5dltlDSNtHcr0K61ExHZVk5gpF2d+J+0d43WQY0yjs252jsLLOZYQ6lajBy5ULQEGNHucZ+yW
brPDj6qd1iKFJtSf/YMLHatYXbvqGgEztvLThzWrknR2Z5VZ08PbbHR1S97DFZb4wM7axsIVpFhI
3Ijt/FgxrIu7nt+G/Q4Rz5nrvgLITAOPMqOwMcvGGO+nr6SlqZLTxZ/4pe6q+S3FpmAVV4C9ERj1
Oqzkht6a8n4pL+7wBcpgqeGq0N/6NFlB07kOlHJdVeNvn3eDjEfaaU3w/3vUrm7CZ5iCowqnMlLK
3Q/C0X2oUBG5KnGuwuyVq/lZlKxUQYnsy/UHGNtPlKypokuIllfTtPMSevFQII4VLloysyhEocM8
Kv2dlW0+69hAv7VE0/KeVtkTmFDXvMzIyQty1jCQLYau3QspW12lS2KeiU3nkUY/8oTNSf2vhs+1
71d6wQ04keCO45Zz66FhS48MRI9fBYKvmPHZxsmYI9KvpqDb+VD42kySTmSyLQUUxLTRKqZTvwGH
9k4Qu/B4Eiu9hTxutiiy6w2zRP0G2+bZMw7tAZldQFrocs3wVtIrc1rvu0nqKphL1XLc2+nzX18y
n8WONu2OXq/6nROQbjsttFFmLxsivenUgHlGpfEzx5h9m53nV7ufEsT6nZWznkycQw1+h6aZvKKl
tFe+pDeZMGNMXUoJqoeddIOiXRc41zKafG4UMyHie15W1Frdy2bEsZS4bkZBeJ/4twpTdPvxL2aJ
Yphujd+NP51FXuQeM5SEWDekwKJEXp0GxWLIxLNzpNhppC962Pow129YL5omEs8gdS50bveadDXz
zllhgNA/X2+51UjHEatSPfSknW2/QDtcfQo+GMo+r2DaK4M1/kh/Siwh7Hbqa6NsJ/ZZOG6Xs8II
yr/0naevtCjl/1PB2WCt9FYIoLsDjN8AcuyOCXRFtzfY7bRnXh3KsQ9kcgxXI1QApx38sPmQLnQD
ZATnodv0lQsKkLJVFkjafxUlgvKrmZEmQX0fMMJ5hhXUSzE7sQbkY1d3oF3KtSp9/xGCYjZcF9Js
E8dUmEQwp0SMDYaM105gdPYcPmhHa1E6MxYp9Hij/f83/5KFAb9cKhdqh+SyAkyXJsNOMPxrvL88
s8P3URbFhhSVJqsmRgztY2cxF3b2AukcSivA+ziF3MARIoRc269hUU5qyiaaUklKQC8SnSzPBjcH
KzL6MUPdXACBPw4ngpTBJFAjEFs9vhEyWuJsaheH4sBskryEz22TNocsSs8IAV+77+iUWeX3CCH7
/CXe6jC6/VAoYiIO4TbwsTGfnRZrBypzVb/RP44XAIMFzDuR8yebBfhL/OIdhWcsxPawHmpW/y5/
Xv0SOO89XgODHaQ5S6OngnTsyeZmoqJUyfyEKmDH5QKmwhq0YnVaDbyXFuoJJQeomTCW9LrQhpU2
D8in8cMhMI3IzeZL/XmvXUVAZiQFc+qUO50pf5xdGKZ0evRJMTFFLgL5dRfNeDA88xn6bLxOOLCP
Yv+ZK8ZtgWL9qqK3TbezDSQadr2qA5JeHoIyBc+3smhdPkY0bzw510HEFCzavo1wTztsUIr/N2cE
NLAa8OVSse0QmZDfeDi3CEn7rG0FAurIROBRw11oagOv7P1SQeaP5SijJa3e5irX2K48jjjl7vSb
2ZYtwWxLJZdqnkwivxeG+tIAHiVe9tgCxNslxoCWl0JGXOGijmMIFNSBzDNB5wrYPNgD/sn6Hk/N
OexufQV8IrgODTD4qh/mt/H0PHY+39JlUFoX9Z4FphcPfUR5To25Ea2rbDzWz7koYuWe3XDvjaal
JkRfXkjV5OzyA1Snxct0Xdg2XMT67a9j6iWJiurGB6ng/+GFhb7JSotpL5wFeFqbn4+6ULNLqJOf
ZjHyyJ3Tk7q4YEg5lJlhh79NE3GRyBXLda95V+yxdCMVY6wqI7U7rHbA2SH4Z/7Y6pKq2gAMFgth
yt+HKe0xQ8uafbxqA01mN08HdvW4Sr4/+d1+C+UImUDqTpecPQ8Ev6uVrlVLWqTzUNfOPtc1F1Cd
f8tcqp82dtvfLOSRDdSUVLMbZBqBUccqlh3cD9B3c8FceFHUMI45Sp72cR5rpi0ZVRwq9e/bN9J1
r72COdZyZqetFvnqg/fORVeTMCTHjE6DmuaG2w6/FjbjJo7dqrsxz/DPQNXeZnvUbM4S95cJTtQu
YfIkirBek4NL9YDn2Kg2mMxgPUXzVTidAF54l1zWOekzzSy44pKH42HisDvuA1pktgfXfUNsQ8LH
a5S2pK2ARCirzUCLUmI3GBGjMMh4j5T74fOkqHReYb+PCCY+LBLTApGREZV72IQyMURJzyYFBHt9
g1n0KaOo4+Husf9sW5bosO2elRx25omAW0+V7ql3pOX65a3JakMcEDRJHoRNsVgzEUWhfaRQ96Ya
dyGSSP3R2h/2sAGaTM8t3cfk51yvqfY83bpepLuoJPlf7iTvmUYBwitkrf9yOyMxBMVzIcq2mJ2I
UMVOhIW+N34WtY5IELYNcF19ixBESyXCYjm+mhXRUcCqGCNqXKDnp1H22ZZw2dI3wNqanRoTy7LL
x0n3TbMl/CIcYV1kyL2hPFc4qKBU3pesW9pzQBY2i6GlKhodPWnWZ+1o+tjVFPbz8VUm0Xl4sLGR
H544MLr2tBkqAUbFQ3p3H1Hd1uwLyyFv4/OmT/dMcU9KELfLozW2bnsvOWVGchaBEa4EiHq640Z3
67LCmV6O5YfdUczQxOMhdD3G2Ruo70A9d6+LOnZ75bFVKTJ35rNmUBTulKank/Lg1crJBm+6mPD5
+/6vB7G8EkO7W5h09a/zAq1rBDzCfeOB7qt9uCtafpyYpiiu7PozidmB1b4oKHYRBF2MNOJRU35q
MDRCofWDkdhCzWzDVt4qaEYcOy8zVP3O5sbhaP9OostJtwjuyr+STUb7Y1fU1uyGd99vrOHr1da8
2Hz0klMkJRIv1043AQ8jJBL/VyTzWmKQyPtUlriwfTyjbxLq93auMGBCOIjhVouz4IEizNB0Jm8n
1ejrNoeX0rfOFdDmDPU/YxkvLX6dkDFfRpT/M/NR5L6qZ8FWBCTcofvCe1bW15NTTV9aXwOWcrK4
3Mjh1Ch6Dqi40K1ROeiIaus4HGDS5/GR9V1U2XiPo0k5Zn2xLiwJ0fhnIpZWdA8qgpuEEXEEVN9v
rMFTw+9vmsnbOzA3zp/vUGbnbgcvQSZ9tYCOuUKJLLI73lkla6/QruwDcFOMuLmutoOCuO1KCDxg
AmKebAncaycIalK1ygA+zU2/LyPHMCRTS6d93QOOwl38VY89CW2xZqwcfdfrzC78jWm1noJBoWkO
y7Q43v0E6F/+CVpN1yynfTowz3+quCwvMoh0xEicI95ZAEE1iePkO1S7inKDF4m4fUYIAmg7iL9S
+nfCvzahh4/Vw1NrUrpO//MnDwo8cTsLQkLBX24t39K1w6x2Mu6GRqHpd7rBGdZsIb0wTb9sr3fZ
Uy0LcqzTO6kS/hiwEqMFs8LlYt6zx2IQTyGserLxzMr6baIF9nRgZ/75b3Hb5B2NLr8KewPccE6d
9yMGQ9i+7nRFjbAQdGBbhVSKmRm+QKaLZ2Odg1ufN1rKKAjpr3f4AI7FwbPN5KMsAyf2uYpuuVPi
hUSALAQepUJEAAWRc95yx5mmWKhoRF1i4pZly6vDAi3wpwVDsBTyFdxl0HBcH4mfTCOI5obY0fMj
BUg13h5x3abrHHiAiZHWeKfAqgUKXEEDVAe9PM22X0J3NCqK7zcQ5+tsRusHmye7sARzy0PlTQtb
q+v9S8QxXEE0RdrrU0Zn2b7jRy2IAnJW2yHaMwPfRzTytnWm1okgOvp8nTqWimhmocTwFh74XGtZ
pudckTL9jg6T/eZY7iapw3wyPpxdaUDudqThCXApCfBf3QHaqIWhjiaeZDTTwAYL0Va4+71UWJEp
A9e0Q0/r0mtECs3pnDeWW+JaNtsZZqhCsZ1ItC3/RGAB1IjFhsJjnJuqloJJU2CWDMYMLC6KjdpN
MZ8Vchxc7427TghHB1WHVmRHUTNiYx2MfrD023LtzV7ujFTT1W/M40Ltkm8jvp7HnFNYiBbRPtf3
SawUeUMBS/HEtsymeE/ibK4hYJz79opO5SkzYxM7Wx0hmShMpFizdRi4L19OlLMoNARFkR2pf309
HAa7qHsyBjaW1TBPWsuk/6yGpdeM2wGdtznNCrn1bH0mhDQ/8Eed6dRpeDYZisOw5BLsGaXq2sNt
FkXX+3q6wX7B3eZbV1NxedhdpZkjPrkcrjhRfMhppy5xCUXtZb+ff4xOr3nM/aMjGjgC3Fqi/qNM
15t9S3gZHuoGvKYffE3S85gn6pbUw598Xx3DVLuqBqpkxA/oaec3a3MxgxZID6DnEVwpPrpTMHYu
IXVA7JA0PrCzw/cvYiZBmwhDt8F6SIcwt9HEjjAKaMYkiHdo2XMiRwr5jf2SpczwWfSJojWn6hFZ
Y+Gnj9IFcWwx/c6NU3C1vecIQVNHL50CoTO1mB0e7WRq+dpkJ+5zk5PEfb0huKbTCFVo9IyBjrxl
WZDaMYzU4zLVgZkAzmRV1ICGEyH+TMuvpq7JEqaYrzqP7J/H0qQlp7iLs4xUzky4kqI/fK/fKph2
LVWk0AvI+7f9z6RaszwOAYf6KI5vNeMn6jI56fv3lLvqIvKvUZ/iMGMYt1OcJw08uQvC+r6qYlNV
L9yQ+Bf70dk5A6GQxzsKO8vpXjkjVUCPEKIvokiC8ZJdqvcMjXTA3XBXH80W1qKNpjuz5LXFfy2t
bXRabSSCoRu3FBurYqyAQX/PdU92/HV4hP+zUX3Ls147WxuOR9wjefkDZrONclWApYK8qe+HdlR4
B5Cdk5eJONu6Ycq6DV2u96Y/1mBTD/GDPvq4E+5Eiv2V0ezRCyfnSS3UGQ3m9VGD19e06h9wucxR
sbs9MqWiAdQ3Hcus8rdX/+8nozxIGhk2qiaYKNBIteS8JpAXJ5z7aPuwo9s9sdqzNTd2qfFYIKUo
q4enywEX0gZInrUTprxfAdDox3yPJ6BNJr4PwDYSrLIEnIjY0VHB9xWETQUAGfQpwy0YgtVY1i4t
QraQvKFrt4VNJclpM/rlXmyKKVVUIfgb7WyfCtTIm4ZfSi4rutab84NHRv85GwgFwClSoJMEc2/b
U0tesHrBkz62evjkNRkWpbMoh9Twz5Yu0O1vXrDLrkSGCAa5eVg23uibcIF7UCiIFR4OkVGRWQJU
7Sh7b71gtU5sez0PvQYlReNI7p032A1H6EE34soueqnrAacUPlNed5GPl+hwo5viWTSzaEBveOFU
4sI3epUjDuMA3y2NI4x+sHen66jfS7MK9lhznumc5yeqaY7V4mfvxHOHGPJ8ZbKHRI57n1RF5kuw
47XiaBDwDvgjAj8U3ayy3gYK+j0xVgeKLzb3Fv+9HHFJ5bwLbnKAtGxtaPMYtultWVkm39HNZ2MY
sVkfvncylA6QKDfaiu/3FUi9jpS/xfSHsssLAx3LokeZNQE+wzGZf47VhTEqV4PexQRTyUmQVvQl
WdrhDfgxRSHQ2O1IHw4DwwqvJuF8+UvbOJ+OspHZ3U9l++aJoOKhWwL5ACFlyWu0liu/9TTZZOr6
1a6cQmhqCxjmdj0fWIa8SYxZlkZmdFZG/K7qUf0AT1fKgUY6SpFUJ86pqg2Z/YpFyTO8EoihBbI2
31nsz8WsDvLp4gTKoPyro5BDagN+uDAGmuYvkktymqt8QfooDs1LIRYXKtaMDsJdCGWXKTHX6cMT
ohZV6pstFScbUInFunxEwemlm4s5o0Akg8wrraVlTZvJhg1KqeagliUQewROQeVl6Ln17p/kOWe8
KLj7UKp1mQWokh0+VrSSEyAcg1lb+Sb9/q8V+WFRoOXdOnKa/As8BmKqTK2XRR2Mgy25yUIntnLb
kngW8Fq/4u7ncBMuPhJhZaInPM9Z0udnDc6KEFeTjv5057MtAeYKrRx3g/QGPTEEkjTGDrmFc51R
rwd5IVdyumZ37zLhckXgIvTXenEHFM4NNEwf+TBT5KkV2u2iQeV5bXt199o6iQIpez6LjST96iNx
TNlho0r7YgFv11KrYgRWG4qnzf1JTnybxZ5WHP6BeowWS2z0AEtDpvLM8wUjGOmF0uLHxneonU+a
HBtp1c/NN6W+tVzypADCr/Xs8q4ScPvfgoekUfnUjzmNowISoh+AXIaudGD2Ij+O8Gdj+SRf/doz
89I3cAigyNs8K6kKu0WPjmumB0CEwEZ4Cff+MtSDZ3gknLR5Elv9eHWxef3ysYslbTj/nEqcHRKK
1tTNq5uE4QAtzRYOyNBtwgiUQiW2nSIXIczjKR7GQMropRGII3HIxlbzUYVbDyxvBFBDCx/rj3F7
Sn8AImCMsWvZyC0hNVMKPgdG863KaoErLBxi1JzwcgASqj79T/lUFXvZypaV647+fT4ff/FkKyjL
WPKWSS2V0JoIk9GH/f0heJ6df+xomzUjJOnzUiHpOiYPwlKFgvSYuVMS+jw9sp9C4pku4hdTcZD0
WtXIfWZfyGZgCUzn9gorDlJOAVu4jneOgLYcHlnPIhnAiUuwv8Ff/ln9DSwazZ6q9W4Z1M4+de7h
jj7MBCv8KwP66Y0BwMmA4Ixxtp5Wi5psDkIOaQv0J/mP+kg/r3Ln34NTZV56uHQ5Aq420Qt26GWT
6zEVlPoU7j5eDArPBTQjPQCfo9SKe4DT29rC0uGkr4cB8RX1fDN59uvpv7R91+iLqX2HcDbH28qo
nLnCiZhJzCqKiUAlJ1UDi2pnKs1PJrYVLrNM7U4Q1lNs6ASBYy8BPd1Xnt5WTvZ36eHsN263ZzZB
YsmBX9aRTeLWrtYP8LbcIcirXQHA26n/iNUZYW8JI1nAZ393Jbx83S9QAW+FA1QwT+a0VeqrLgln
XlyghmQ+JQ2Y7nILjA66y0RiteWdC2qivhY+N8LUNhhyXL5PiyReEiISN4WHZaXSv+33kIyiMDHp
T9HpduSiSPrMgvVIhtSlmAy1LTvJ299bd2iT13lrwTV8zgR/OYegvuYv6MLYmNOgjvC7ugzRQAQp
dheil9o+/w+/6997gXGsyfnrMPWHzk5Hql2OHWNfw8nH3OOnZxkMcwgdeMuSSGUEOiykt4rR5vnp
dTIgAYM2t8aOdGQnBhrbWn5sG61o0kvarncfsgfvjoYR7sNSWSQXCVHfdViTu/+XvZv6wzaLUifp
fmhgNNLZtyYv0tJisF/Z0oTmplzWfdlNo8rYzyZcnFhBS4yfFj/5TN4EEC+At13EGFBCfpThUahE
VqaB7jEekNEUrYlfhmaFLY9Ehi+F7cmEQ7Rq5k/fM/Cg8tsM2ebPMvhyglm1JUbNJthaHR2vZd0N
itqAWTLBob6+MZHVaQ+QXqFamDrYY65/APDmDf1sAcPh3hghT8x5CdT/QNaRk4frP2cvh5hsbVhq
Pw+NFDA/1prqNbfizJZrEcJUsjAZuERYjoE4StJQW5l6yFM3LdPjtq23wYwxcEgrEGloRRiZ0jfX
eeepCr/OLbb/52iDCvAx63PlJo2A1SYFSq+U38s/CSgil5sUnrvGa/bPO3MVhYjK81BwQA93z15T
Nl4B4e9jKfFdUW3E/tvOm6OssIgOYggKlVbwqgcujGSv2iz386z9en501SnHpusDZoHGyxzUWqLd
OuzzHYRJDUlhtfX2Kx126PlCGRjcb3RHQckkzVptY3hfKFTLoQr3mwaAEpyQKpgOTElAzhShCacO
2j1SH8ATqA5mcR/O57xRI+KT9aVaTexh7igQWq9nEi6JtQmFEdCdrs0zcKXg+yw4IDbFZ5z7B+f5
Hl2NrsbO2jAc4mPcn0M5yOo/3tNyX/QJLVoG8QGjqlUbyCZ0WvseUIurTxB8qiXGSB8FLBrCaE0I
8VaVev8kgJiXUO3diGhqz4lCW7/yjAtpofwjio3r/H8opfW/BWiJDrQxy7Nx4FA+Ot1Fk7Vn6axs
N7DpB6R2DeqFYgfXGRlgaCvD61LJZ6VZyYnA+2J6o2e7uhWROhhYxSwqOjylI30uFJ4lhN2VzYWG
9ImCTbksClZOlOaHFcaIXHrh6ORQtFjeAkG3o0AbRzyErv2Hvjc+Oqq0Cmv7JNDNQLba7VywV4Ai
WCxVn1GsSTVRp4aI+kVAGdQxN9cJ1C98HC+XZ4IKdX092HraHdY96igJfrSnMrZvzBNw7qI8Prj3
ZTl9o2Sg5gjC4JJvdWN/9GMKGI1pwfbyesUogA0R/hyHUzvpgQSESNMSg5heqe6CrcT4e1X6yMn2
af+gsQ0gpLktOEc3zPbinSyoAz/RlcrTYyj/XilGyCfkDUAzBPf7ToHiEPPf8bJOnQsLl/4B4zqA
mJVDxqw5K67kkkax2Gf7edf8gb45rfZMmD7T5/oUpTVLGQQSyj9oC+tghLVs2VPSoYw8gjfVW9Pm
OL8IoLGqwfC+2ZywvLTe+PTCTSyz5qcXx8MswqMl9JRe8itfC6SDo4rhi3TCJCMcNNaI+c9q6Tn3
5/ZRHFILchFtTZbDuLPN3lVpobkRcd974SCkNCu4t95+r+e/BaMcHKOQnufG0PtmpOjxZ22gtRgJ
g/uPgFj/VcKJfoJR9lfWDH7ItunArPtT/v/XbIkzNPAKJPMFC40iGnVBFRMKwBUwlevB6/CPAGxq
zGO43aDSSclVFu4pII7+qrQFEQjiLiDJY+Fvp1wV3tRmZbgqo26gIWtehaSinxujki9BxdIOFIwO
NLZ5QL/Yf02R9i0mI/90M6AaTSMOYXNkgTMFKXuUySEGVYsFNkavzwtNMIPqqbIVSKW57y4l5tE6
76i9LGuT7rrdYDVrHSxQALjVKEzHBjjUT+ob+YXPbJxw3lRRH7b99ePAIg35VvRGJzQpoassbaR6
9k1P7VCf7Vmyt81nt0bma8xH5Gx6Wd7C8vzdclz9RRMsqnsKQAXUMxyC6EaFGQhKaQqfq2FpnUqK
7nFi3SmhS6Agji7WvJET3jqPLa0gTHEs+xToqS8MaBxuXy4F5syB1UYv98t73fmocoR2EkROM8W+
QVrZZKm+1C4WomHH6MkQR0szIv3UVnWOvBHXXCk3uM8S7JNmAINbOfX4nly98LvRv1J3T69/FaIp
aGUU1s/pAMJIj5AY2b+Yiii4X+kwwwDqwXR4JR1Huo+tNEr4xiv81SWBq+2ypu+k8qPjd/NDxiu3
5xWKgXLGdifveuFmowd5hVZaFEcOh/V0noH5e2u5idp4tqAOIB7ABz4f7boeQTocvPB7Wn9Vn2UP
OvyyjkmrYgsMm9qYgl8S047jTBIg4vwln3OBbMM/JOek5XUFjWo2jUuO4cS1tRYxSU2FXHvxy2ff
mulqLEobMK1ohWinZEBNFd8OhCz0nQNkuc/WOCx4IpLTtUEQgQtAtND0mWqC5zCaPCli0E86mkmD
cxOoj17x7K/yHNpICITrqAzOiEfyr+6ASma2O5wyBH6YvBCVpBM3QASvOtwExM0HXi3CIPh1Jq8j
UMjo2klEfYbd0uFI1zcwLZAaWoLH9U3ZUiUBCpppMzBPu3nY+hOIjEwr6BQ6ThjJLP+OSherKzJJ
mj15dC7LAC/odWoP/8eKHhb5Fm0tv2LwnVWhLNV9sKW29jFQ33+pCuS601V9jRftCfcROvc1mwjn
rmOHFZAFr5JaE9eJatIfeXoEaIvfrmXe0wia0pUK60+Urdeh2ysPxt/4mB2tCUn0xloj+BhqjaWP
jdWAFPfIIMu8w7KWgFvRU5DxWgf9SeH0ixHfliGlIFWBRvgQ/DpirYpU+Ih5tvykTCGffJW1yVfh
/Un9rPFMG2YlPgWJCDAaxKof7I3VXHyi/i4u3MelNWhch6oG3fCFsh/zb3KNKggqzFJIUo70IiyI
mBPyoCm4ZylrDJyHZXiqPAPpvNtzFKcB4JHHOFmECIMkLfL7GhXIHJP0Ip1xR8iobxgiABYgCeJp
J2gRu3bWM1VH8HJkKHBMQbMV4m1URzoAOYmd8x8PIh9qfIWi3d8ZvxP7F+aeCeMch82b2L/aWgxy
1AqWOAlOQfSsUfWH7SYnq/ftFaJ8TSjyfCXHsPFOcLqEagvRlSA2HtRuYXjLFDyvYWRhnlxgu/eo
kRvlAeNIXJts06aXCwLvEAz+Wk/xUr4BoCFBDZHpQLLyqOnEsr4EcgHoNfh6qkjVF7gCkO/RbF2i
FVuo+h9m1fTRrV3EBofq16Sovv8tPnD+se98rd1mw231MN/q663PKZu6RPIpbwuObppQ81BoOXl3
AXYcssxiuDpHRzWCfisois9Z/0Ji2DMMlZTD974g5tssUTVphXzW+i6fSBpxpeuF1gBeo+0gTz52
3WFSqm8Qht8lDajDx9a1p7pPJu6TToOyalOaCSyyKo/PrS0tpDiM2rhPY+JJ0dXfzkaBo3lQ/+ky
mE/0+MJeZ2wuGiQohn4bNJn6wCc4eo1RPIoA1IWbsFSejfY8XyiApruFcU+nwlFwgLbRtkS5zlPH
Vqc9wxQNtjx3i0scuw11okMJKluLrNGdLV3ZBRY9NPnOx1unRiyEwU+l3xZm71P7vZ856liocj9c
JsSZNJZ/8s+atV7fT5AoKLCpAngyKUO4QpJ1jQW/t/p5v20nMJ+Nieb8dMVMlzCr7fY5GAs5Ii/X
ghDMjjDSB51Cc498ppl+3x19ldaYB560r0ofzs/KS4RnldYUgk5tezkytz+zrocJaSz1ScfxqUXE
3Si7eqsvNKOLlRFAotPtqxLTb7rOefcl9SHD3CkGS76n1jJWbtzOSIsEx/TE3r3huQo0YNMs88Vm
TfWlGnR6EmNm66yu4sUgqg6BXiVNc7Bdhi4h5jIb3na6qE9s/CtbxsYY3yvLZW1dK/Oont85jZi/
7E1k23jN0kZBqPfnFw1owTleIhM0suI9xp5VB4HwzQAXUwhbWkjvsLagHmKKguCXTMp4Pa7Kz1gj
qe/fGITobgyU9WP71UvnFKrPZlAOAc6UHWB+LTA51JlCScgqOYLT5ZsbKnMvoeu7RRAn+uPHcXwu
4w0zPxB+3zPK1qqpFrKeLR5vc/mumQYcr3pHSaPMXrU49CVudoIHijHMOMMNgd5lNIl2M7whBk99
RystjYXHvh/In48Bm/xUeo30ARAT6lCgNkPD0HbBZvRyu8Y+pXJKQDupggqLyqCFy/oQNhJbKELI
2ML/dCGefpBcuQsZ93NBicDwYHqxOCo6c4xKYByt7pGmAhBili941RaadNnaEpKpP/mNQt4ZKlN+
vza7wiZALUr4EjMWXqBxwPemHZBPGS6j+Y2rv5XZzcfV6qeIkOItHCiJ/BpeqETwp/h2FOTuiS+P
oM+aLsz+BPe8s4rIxiNTu4Ppr1h0Pr4/mx0gM+pL+KopTU94G7q9K3M500jsR/FnOWBztbC5vyg9
mgOBIp/5TDhMqCksxOAGbRB4uuAflkBvebW22u4U1h/KgVnICl+sXpCkSkDJ+2WNPE1Ipmq5PZ1i
Oy/cf6glX7fp7reNC1N2gp87K9OPLpgT7c8CQ/NBBu79FUXF+Jj50YEukxEoa6nngDXq3PbjPf5a
SH03/351srInIuIxWo98Vss65LiVlGenidhEay11TAOPZeDZUjblOiu9W8/0feJaas05rRUYbaFb
Dh/hKGf/sfiRrmbfrL5KMmLrjma0kqABmrZYU9BGiaZNQbY1+pjLXOE3JsVTCqRyt959n5sF8Ke8
C2ZHnJxKPpk/lUUaCoD1Ua6GJpoBMCj3JWOWNWYV6t6tygFv0VACGEGT0N3LYcQhLUO2Lhg3HbJV
UeyPIcH0WQHlP0mwQRgACTRGiWGD3TA0tjFilI/blB99IMemeuYXOyHBWmDNzKdR10PlXnjcPQtq
KdtyYOYQvTDYbFXYsDigDuQ55Dy6TvHM6oCIfw9wBSZ6JQom2n8f8y1F03y0jDz5OMiregLfchVR
025A/RsY+xk/BnlXBQHdiOhZsz3bj4ntOo7WetptqEx8vEolaAkhYwxdcy1bs4Yn81CxjOMggaSQ
gTcjA6W8irPGGAKU5++ekvMSTFVWbULYwceXTy6Nb0OS7eEnpDnOjU+F2EV/X18MEFZ/BN9/YNpb
/tX78EQpjpEFHjHS+iLoBWyXhZjGiSiCwuoy/uBWCxuxcevh43yyEac/hnOXiQxdJrIZETNn92tn
CwwMVVBOQV0NZvspxGwjVsl+4B48ly/P6Fwlzs4dtBzrTr2re3kiei43LpLPbN2h0knXsqTfr7VG
SLTOx6mJnqJagGp+gi2Y6imd69H2pBrDDZpa6pV4HdR9IWQCZQ4OTLm0oWS77g+hHMYQxse/8k4J
OJd6cCRfvZkHE1kbuoJ4WxyYV7SVfWGrIxG51xhCAUWT7Z4MrSdDChuWJBGIfM3NBwaFdui9D73t
PGs6xrYUtV2k8aa3Uv3aYWTm4vG5tFdv2hehRRoEpyeWgtL1lfK3eSnPEmAlzEMiCHypyd0NQTs9
6NcrwZYvVmXPGGUC3S0wTMyxTKSEnBz9okyE2CL7ypq79qKLJVMtpGZcd1hS8TV6wD6gnUAM8YX5
s44S/ptoKrcxGCXJt0FlPGNtH7bHWyeZs/S0naww2T6lzo8Q2O+zz5wxlrhg3T+mC5sYRy6UrG4Z
eFWLnhSH5M8v82yJaUqNdPMhvDUB5mtWtDi+xhCk+DpmRGZep0Y0YBoyC5U+zyWohS0bvvZun/uE
PSzYylt3ske2NnKp1aA/+7Jf3cY0YgOxi1RQorqcpir9gbnmsZgMNgphgv0y4yWy9Fg8cjefY6FX
nsChXa8s3Jxy5f9MJQolOcJc3gwvKNYOB0fvexGowjAqrmw+gHQI8Z4p4EyUxzNc47Dl7bMKgPXU
tXKb1pyu1DFd4dcA+b83OkfGtzIjgj8n2jQVj4m7rcAUQfbz8yoLz0s2NZ/ioiUg3oUsWW6rU5zJ
cVwufLeBIXtmFu8hwpiiCAk3Uu79cmVZJbhvSPwKKApe54T30QBfzzAGUv3iRf+uKCtq1oTeNtqK
QkrI47mx0CUs1LlHbaVpgNI9HMoLkdVbU+I/Apg8H6cTLI0RNd41Voyte7h4d+H+UvuBMQ9J1uz4
ebQEvUXK+ITUZEeiz9Sq/eXzdiEg9AhiFMrzzrRnKjgc9RTlMvto3RKPnraY5VXuoJhd7OtGMLis
PZeLqMxwO4xR5h7hnxeW1MgLvN546KEFLT/PnDm7fXqMKbg130Pbw0fiQWwIiAxSZ7AEQOcSXyRW
4mAhQD3wvArl66d+vlPnEIl8yY41Ptg8yoinMq8OAkBPov2pfIJN0dHwFwGRUi2Qt/xkpB7TgRTE
dff1xlYS/410lDjLlueBYyekxy6TcgZVebsx4rHBZXPZEQsvXnOKjiLySq70ZMjypaXvMfHhXx0z
hzIrvpO6VTh2rRr/4gCjCSxFMK0iJx/wKj0fh2PZGGWB18MCDOfa3rymMHd04D+eLAugutDsMLU4
AQ2qQ/ItOTzHjJCexZ2sOJlZT9W4IRZRoZKXYdfTDt2wi54brS02U3ZrOVn1mJZoeGmKjgxtnwe5
sz7AyWhllO+etQlBUIqrkQghBZGjLV3OF1ZWtUDXUz7lPkFRmLdNod4+SLcnhjVexWC1Pt6ElGxs
EvLgWNcqZYFgCAhnW+A7f0kH6T1oNYb6wSTGo1YSYCCRGnU6DjQXJ8vrqVQKKineD4hXUd4+JdT3
8hi1YB06Djg8Wl30I35nnLGQZZsQ9DhaH4jiig+pkd/aGSeEVtVpS0nynLXY1bW195DE7bOD/iQx
AVU1dWOvmLVd3MaJ/yxnP9VXI1Z05jIek1tH0p//6v7FFDCJSw2SPVBT31fjNxiRPNlcKYQB0UHe
1PWNGmZtNygr2KrOsLGs1nTf+x/jZel1QuhKFWKmHZobyay4bFk25IJSfeo/PA8KMO1Z1wGqmfeA
xnpwLrjdhdgGLDbeYimNhsAMpJVBAOY0BK6JpJrKt/JEd2ssEbeC3NDosSxyfDAS0keeaEkqzP4p
0WLLc2Zv/IPqi09qqzWHLyIX2QQOJjRsT9nYap7EowSAnFDk4szaAEMAmAIyOF8WYKeN4D/ZE8Cb
fzdBOpBG24ol0MocNLYw6IP0ug2Fxma/VhFe1Hms5ZLH5fSUiH4RrgLhUlanSgyq8dNoLu2MMyJS
1JToZchHrWV2dGs9cu/e8cS457Z6Ad9DI550o6TVS7edxU8+p/glexr8ALDIPjR7UYE+SWBJv1MD
P5PstzLVzDpZrBXHrVocsZjH2ayGRRhr6Rw7fvrnQO68s2hPDjLjXRxl+NznHx4qDPDIwk8mIOzR
tThrpzC5jwxHmBeYh+KRa7xE0rcX/pbPolaaO/kzlMg7Ct0sWPPElHqYYKpBjIlsq2onnPy2iHYL
uFAfWu80hopfBRfEglkQV7j/U7FEcQ9QXbbGl0+J+caK11KPsp+koWM4cJ6pmPf5BgjZVcXyz6lC
KavOSkgdCgrPYMAsn0xu0UG1CWmgfPf8Zz/beyxgYP1aV5k5GMCSytbrW2PkjfZZk2/IdkPDROxV
AzxFHGr6y/BYOiUjyFmsZ6q58k/V/LrFSlsRRxgq5xh2Awla8euMQdh6UFQZBtiVyUYwP8kA6aWS
kuzzKyP+8/nbHt8FIZu23E9CnYuGrzdxhsNF0T3cSe0tmG/5TaPPYpTQ66YTifQqXDDE3dkWicxK
cBZjpYGG5FQSPRSS3IkJ5yG7LRs27l8FvwxZjxb0RmhMm3dYsubiRUKBgtArIawPzaVgpmUcHAF5
J4tXXqt7WmytEEzfnh88SBJqTdRKekIpFt3xe4ZflgZ1j2kyjDZPeQ7MCDL9/FqEgbK6WzP4vipF
+UdzZCRDEMxVGyEPIwovHYyc8V6SwDT6xJLuWRXsg3h9bVvghhxqGCM+MmlfrQX3NqScYeMwcILA
qM/jXml2B5lLszFJE31zAoaHU029EKbsgxO8m9GS0JIOmJetGKL2X6Ym6aWHj0bgmnbCptMAXNay
n1qcIIfVJOn8cfE5MG5N8zJeoYZi3iDXmeZhGTrF6sZbgnq6oVeabRc4nalkuvPY0EmBmzzfmdjx
ALTjag0OaiE8jnbhh/4QkODmpBhn6+PQpZFMLHL1XFUCHGtpOQL898lyNvQu+VWXftRc9Qusq2J2
cP2juTCMjxeYaMviiZAJ+qlb7N9EZ+2p5CsRL4OVJVZbgnGpeeRuC3BOfwviB47Ww4oB7Ozsz5Sh
AKKdMAavZoLd2bJ1xccBVXVazXJ5B0fgOft6ZVwC1rKinWscDBKsg1Ol5PrKNQcXK+YwBDVkkVbw
3ZSY1D5+OnOFkEau8sDhZXV3tMrGsmRKfUpU1/b9K+IugtLQxyywvaD9o5GLwTVmlEy6TRcXllr7
khPRL9x4oqGnHHZRMbXcDpdIv7RxoNZZ4I793+eAtpAQSuXk0Lwxf+GdLdh+nUeHp53VGC2LofLj
RAVtLalD9rhDAoT6bhi/j0P8NlvSZri3CBaXVQtjI2JCdzrfuuLZPWu6tHGEl5RxgVwMu1bVXEMH
nsc4KhyJM1nDWkWZ13FJKwYv+8VfgXI9n4zLVe/+lEcpgLoP4vTiuWwcMA98vy9z0LikxU3xGKgd
P4JqoR/x7Ceboj1zVQOiu0VnMzzxRAiLVnj9vnihGbSUIINrtAkNJX6cpHgT9tETlTH1F+4BxmPr
y17UIq64s8aa3pkujjNlqIbnLz1PgPOMPvdgBQv3ohocJglEwpXZpnbvGWTD3Px4JjRkbrbcJCvM
+rmYdgsesXWB5qcx5oP7fjv9h078aYoZkitAgldutx7RIjBtWiTc/JOX8P9AuA332kOn7LgywV0i
UkX1SRP1N2Mwovs4kLXaibcOrBpZzJUdPio6PHQCWd7rAsy4faa5yDJsfPAU8vUWqzo8Jr4cYhT0
HirAOzKDWe3VuhhP9ONZ/5M6XNUXjkMG/poaFZiOSStmPTtQf7+MfKET+gsCtvQxWenb1lU0oDtt
I3TPT6bMKegmuKSloZVoBYrp6FdzLK80D691v+CQJFZ4KBfv5h6VOJI7+clb/lGfN2C9burNhQz/
Kg5u3q6I3z3A6MexrydCXJSSGBPoshP4cVMpWV2LMqDEnWlvFE5nw3miK9oC5CT9e2/aepQkzq7t
FWsCAwBuRvC7UI7NAS9jhbzEnp6XfRAvgVuMb3VGYXmvWem+kbRk5yE31lhnYiUbrCc44Q1BTN9A
fnbYCFxWPNdSyizUBjsXmWbqn/pokwBXp0I71zA/263cP/xIu9kjqB4dlJyi7mYaf85tHHHKBf1+
RIAoOx3X8QuHCz5p+DvlgLgF4P8p/JZBz7eF+A1nKATvoS/pAMtsu8fDJSL1ITXNGFtKQ2B5v1W0
rFU6fsmySeen3aZMuA2gF2Krpa2CnJDXCQBiju8iw/GGoi0z8A2OUsLrWdqoS+5E7rJc8EemCOfZ
Lfum3z3OR60biD3CVm2sAIz3EkO876bVHMtcjNJQengH23PFQ09me8rEd+eRJakw2AkBjvZ8jl7O
qLR6Z2TSYwaVMihpWw7DImIOyRfB5d1iZQ/JObCw0sIXyEPU1xezE66EFeiM/CStZhkQ4GlCu+qy
0eN1/lWplHHUJ8gjkXtHRdzNv2B12dNSNngIs5//kmd/qlGwvq+Kw+M3cKAle6nZMP1976vec5zB
xddcmlkMEbxg+eTRUTZcKEQ/xtrG8/WzKxCdqC96YWu8Bv9dMzkmQb1A3rKkKzuGNIxUCTzu9UL+
aoxprfzqkPU+BsFG23OqSy/8WJD4VCFmF4YAR9NBKz66dOum4OjvvAYInqMAMDbfnaOpK7Orz2eQ
E80Q8ciVORkZr+s0qqVG/sYGpuOwk+Pj8gdL+0HudTcMhTN2601Nt2jKckYLkO5/c/LTKVU6Eb56
nkDuIp3cEeFO+rSrmuOcuaKo4BUjEyRoOb/S+kRqkUjZOe0c/xUMbvKlvhrQEDEMNS+GIJtd33rF
RySONJZoKu8KMcQYp18usPdUvk3/gaG4YIyotbqfukKgd9vQEsrwQUIdhImEelczrxAeq+ELvqBQ
VO+W3B+WQOxMdws+ZPC8+oywSs9fVibh3nVOd1R2j45uLPlY82F2+nASNbnpu9uG2SaGi0Ln/Mwj
DQDG+dQ3w005FWEcAng2tE/iWVI+IsoOAUNMRG6vdjZMiIF5LpakZ6pLXkBMO4bu3U/7ZLQ6X5qA
Yzhf/djom3auowB4dRBAYKTodbahipQzGVm35uBdyZPDUyiJIaC66BqEwhLf+dnRZgUD6LYGf3QD
8WsP0j1F7KrOgqztZzmt12VOs9D+wSyy2Yo8C6u9+/HYCIDw8LA9C2iMK/XLVvxrSujEfmzkOHSR
NUi2DCJX8j/GoHgHVAZNcTuCYySXIAc+mWIdF6yeLZqGUKL2Ghl7VYz8QViTIwDKJCJLi9RsflC0
4JnATi3WwhZXdBFNOsFS5/MkyA2D2vLIC+0YvJSINx+g1/vAodkeUg8ENW7LDo84KGwFmh5CUeOS
NeR4V6XD7+2CulgPD3yMklh3HFDM+kUC9BpLzlwYRKdc93be/C6XY9TizMf9miYhs6UtRAXVOL1b
kp7978H0zkZcqM1anrAwEFtGi62FC0Jkd7pHT+rlWpAfV3ruQFHlXKYupaxsy31hfmhhcl53gNvA
tRdGTtbeXvZlafyPJtO6YiiWUPOkUqNsZkVhF7+prmsa52B19zuKBzxFQg6zwej+vWeKtOKelID/
ZWb6l3SFAG5OzRsk8a+1TDn7BjyyMUtUa+9wVnkx01EZetRX5UbvFRftwzMgemjtmg6k3znE/OML
qwNgie3x4wmOLANEVAPe8k1Oym4RB7ZOzJEhjozqmZQojDCvj6dfV/SMBQr/32buB0rTiqIaAXw7
Qg6VU3ENVITpaPIBX8a6k5mntsSsGRwHSfMY/9olWuggqnffNV7MLH09qUwTfuPntz6H3guLVByZ
03IfzMcNLqDFrBVYWRkzBFQv4guAp7IaQWDR4kd968tmxuV/d9E9NvhZL9gDGV4V3qdt6cfIHwif
SiZ2hTRmzE+JtegkDz8OmMWoiA45xLsuLr0Ecuwh43xQVfIdEY2JVHHLhaejS9JRyiLBr1aHeW7i
tW/1v1oZES3h8DhefaPBpOE3BjOjA8XJWnLDAGUqreKfo4qpQsn3f9X5TaHEGdyZLQCWGD0rfPRQ
NSJE0hUSpNxOLPrLWRG3JiNg2gvsdegH1WX0AnQbf/z0oNcY6KWvN15o89yY4Tvmp9EVVYUejHmd
BTRAM2VsWU6oVYrgBJ8hzz141RtYR7Yo6xwMQ4VP9talRcAFJyKjqlAl2spGJ3+nQzrXm8JYRc8P
SEUXZXctdStmEBrhFmdGjA4cOcbjSZsjJoZfK1j6zj4Vyvh7DQsTogmn3KR77DFcxNuesS3f9zDD
Mp0Iif30zBE43MXFwxQep7QI1Rn7zWIgvwnlRXcDY4WgfdC4cswXs1Mtz9iDuzLa1fMWDsoKePVo
MviWlzDDOxB6ljPV7sTkztZngYX3kNphINrKUJcvHNXBVWmL+v9GxyCnDiX+nmrICVSQ8gIJIz5k
GeFtwU6cvg1CAQvuUMf8BvCE9ME0i89KQJTepkcobvc4dTZd60Yxa++VKUwtDGqTMGRzo3cVOffO
s22vX4IR9N73orsKaZUeJ7cgx0STmLNiNfTjMQmEgHRd+pCKjSVJEGzVK2ZblTV7xtdpimXvQH0A
NZHtG7UR0rtsZ4RQx6w6NCwPwaCR24pP/Nvp3RtK5m3jhPRP9+SUc4KO44aBxnI1Y86hwOrmxgTq
1uU6+s3ytbnnW+bPL4h73Vev0wXakhj8bLlw1I8LBZxB2heh0Gv9LUKCIkdfy9SIm7g7B20r1/ws
unRwM4HTilnyh6XRvjHmRXcYtri+g6gGLOOLwwA4hcQVo9GHuSdtCMG3nlgbaVwwr9iHcAX2fVNl
hN7CT61Vhfi+BShzshgHu9vPfUhncayuX+Vxl3vsKj8M6n4zu+OC0FMTfMBAayYAG+2IWZhjyCnU
wf/Mw3/KHBOicpBCT3uj0BSl+q73vSO4cxvj8LNoQ71+xBzdEcw90Zx3W3dL7MSdq5OpPsB8UZNr
vBi7M+vtb46oH266wxHxX/3bM6tgetgZhqX0mlAaYlQGIiZXUYyCgQGKL/fQguB0oH+UDkmnHTeF
DD/YE0YW57Uz14DBUCEoBj2qnGK/bdgCXQofWThGPByZFdgdc76WlnHa8w1D4mXePT5i3Dh8r7MB
6yFPRjta6uQNhpo3j0dhKC6Jke4eCscsQe7eZSkku6XBVw5yl3mUN9xeLxbTSq3dbghDIYCqeJnY
MWq0omsdmQx/ob/5TepfBV6nItpczJai6ZZgAvkPzCLPP6WVxCghvaMdphQ1QkNMezaechS5Fz0/
EMNGwjg8BO9Y5qVIyg27s7QHMdw/ROtvZATlXTXVvprZAlN9YK3I3toalNVhAYAIu6kHEHIHSDqO
3AqAJpOUqlqwtpFkiGO0b2tUb9qCsPt08vgpXAyDF1+WH04B95tk0OwoLolC/zTGaorUcvmz+bK5
Z1YynICR2aXBdVluvcQBJd0U7/CdEKH6y2Yn5be3BpSL3hdd1t2kjFoIqQta1ceVvEGgpShkpzpx
IyNvESUlE0bKRkh5mdJm1RLmpFiCDrnh73nsNd6dVkg7p1Es/R3lNJ2t6rUaQK7f31VqLR1GxZ9/
HrQrgtaFWY/T3MmpX5yMJHBEvLkBlv0UQBQx3ye2dI+YdSqeA+I0y5bk/QJsX7ldGbP9+4wSAgbO
fvSXU2ZjDrqn0OM4tTltf942B7numPJjxzitzFoYWi2icCwHi4oekwADfPgUZUwFB/jswDH3YZrk
kkOAAxcX7fVC8l+mQV5DsYkwbZHM0+rn0ZJsMJkEzM0fKzY/ypdlcCm+cfkmGHUDC49PK4h69pBY
of3vAIKEoxjLCYxuJXCMEPQu7CZijzRz11tkChkFn8c94FYTgjq2+oAxxHpkoBiI4sThEnVOs+Xe
CJ6RLXOMuHsBEI34hVCYFPboTbCsf7FSNJz4r67NpzSt7/6HbRmmKVurOEhNbllo54A6zmF1+tRD
AAK9noCL35Lgf3i9oyaNKRVjIfY0se1LN2agPVy07b223BzKT+6KZoPGlUjA/vjWOGYQKoxpgy5C
qpRW6z0N2tDxtoacjqoA9qnD1QOHVOmH4FFw0MeVftaWLq4zjNvTHnba2ejOeCf80quD4sBG/STt
QyYDLw3h0FvM/DBH0QhAAsjp6+9xAPkajbqgEFfEfh9ylruGHAvraY0h7gjUBJR2Ucy3BUU1rHOv
rooNEv80+ij82Ygw6rNWRUEU8U77pXAY9P/W9YFrNTRHFP0ZoWbToG216006AfkBNf7st67OwGQE
G2+kwL2l0FMEuRODvB3aRbjdRu8nrQt7aq7M3pgO7TEm/pTfbJBxMDyfoqs9kWr7BcZozIqA+27z
NhP9BlnvgE+hpF75lfQ8g61k+XaKbFjnxRE4vad3oA0MSmDAS/V3ejds2Hicsyjx/VSHDfOspWz3
Jhomss6/AzVB9w0PK/4UrF9Ad9dMLjUmzs0ZOV6v+TmObWOAegEEeF6U4xGgnGPHE9b4QQ+xvKxN
AVu/VyUldULmJwzLxfoE71eTPwy/Y32TRcux/6eJiOuUWysJuRpSJPbSqy+VPWkNWyhy+DpJzbHw
wRSR/XZjeXnPz0CEctggcoHHgunveVMJMF6Ryv74ZWdpGvWz8LvUOqEaGmXhjFJNHSRxWW2MgdTw
0iYbI5gTt24vXigNvNEhMIZ3DQl7yoiKMFTWtP5ncCJUsIy/IjqQucPxjVq0jRbhFhoT70lkKnPT
CPglDBmj/++sjeilWf07SqcN2ydA4oGLz+eZkZ/HbYcSCm+KJ2rvQL712vU6k9wIghxqfTxe2QNH
c30qZg1njpB7oe+cgfWhPAFGyuUsr1GprOOWV8gIJQAWjX3OGLRNeufcdygrhkfulbHXhO/k/7Qp
pkdkGziVkWS5RpM48oWFd94OJ//Qf0zxa+wfQ4B5dLwFxEB0aeZz+t+9FijtFvO7daxJPwxCTwgt
BWx50LOSimQlttssUUCg6/aeTG7iF81grbdMegANJTmMdUHMsnjjNn+YO9HBaIpUI2xiSORG7d1q
3Q5/RiltvuTnLBKsU6MdaSe7MRhpERiBho+tnuMALXZnSGYUFKDwqbVF3S4QFGq/jDXQYD+D3/Lf
MgmdWfOVcKPzaHKct+HFAyYDcVWtCXjiWOb7sjhVxnBvXj1rzsqYR0SnxaZ0gLafIR5WSIe8wnIt
oW+fwzGbpxMGHFs2RFtC4bqvNfmaqL/agWJm25DT/T/Cw3t3uihQWPrwfsoARBmcCF3+i/cUUxSo
lbKxqyOEiVhoV5bROhY2a8AvLsFBV8mjKL9Ba667kwt+rh8TkyfH+j6U2iR4sBrDE4fAP6ZIXK0I
FamZ13BrjypUm/q+R+RiHe0cC8Bc5cu5U/lKdCHBWMwzSDsEY2/KAt1gTHrFwQgGEhrfU0BYKGny
wlskt/bdwRaB5+rkr9XTAPLK6xaCjmIMcPKovBND3EoMydVi2bGRNAqIbfI+roP0UfPZn5jCIo4z
CvL5ib7BmE2koeD5T5TW9vz5Siodw0luSwRXPzaYse4TdUEaN9r0fXiwSPrIsgQbjPOlCMWc2wKx
K8V7/quf6ZVE05dNPXfxPovQVAFbarC3PJe5hR2MEK8nuO0fxmHJ1WHVad8w0j5kcdQfkMOvVo+1
hXmuojpCQU9+mJ+pIzXHdKsG27Ol0W10qfWKpEblutQhrZ2dQWrWyyzhUIfI2lLZaIYV9bw1lvxf
kxn0h0HBViXPjSKlUqCYgQDsp4QNJKv2v4wiMM18AqzLz9B9mcYdl6K5634axnDrTkaJpkt3Fl5y
rpaSCd5/D8s9vMrvSGsEn1yFe0/5gvlQPE0p+PK51BylRtwOcdtte3RdCOAeFA3YOcTqri8mncMl
7hSzyG42u0zUSrOJASXqozPj/KcPrnFtxhnrsaYCNfaNOw5r3HmIQmSIC/2IVKBAQCeU7BhGlkoM
E/HeClAiwCSzMzK2dTN9L1VBOD2f9XdbYZXPC/jdsoMoKjRh+gJDMm1zM2HhFWauBuZI00+T7k2L
q/L38b/77YGdM9+ImywsNcXFNjOO+Ikt2U/OgMUBL1O5zXTmIWZsG9ChP59dH+c2uNPAdEsA5w4F
e+uAPHVyJWEqfhm+iyzNiAq6xpBUlkt6DGLj4cBH2HyJxilSxrdQV9jAPPzWqXtyMrkRZ1C0CJbO
CMNMox6uPCjg+0v+gy7c4wdtWeL3Ns4uZgDLfuUheG8s+NF5AEMj1kfLBCsQQOj+Q7qGnxgO9so3
oTimH2idkt72TM9bnQlNrNQXU0XCVCjRHiCoRuPFAiIUmfdSM69I1knDh8Z3BWcHRo2BhkExPESl
7J0gmM7LHsSLjUCTp9EOfmFGWqh5QA5TGdS3OR0eF8heJE+80OxLq4XPHL7uFVm2Hu7A+Lkq/QI8
2fM7ouE+3WL232guA9KMFFCqwOSJTd7Fs0hPzsMnBec+pLbWi9WtcrYuZCXq15mNu5hYpopK86/i
kEXWd1p3AJGV9uodaQqShxiovmZ5tLAHStiA9UVjrYRU/vzxGGAI55yE+X8uWd14besQT+kAe5HZ
iu/hQSVwy92xJEq6UYw+EVsYmTEe6EyL1uT0Nax0sAISZNzJA7fC7WYgMulYQjREX6rAX9ckXvIM
VW75XEpZKKmurIpZZ1PmEuS3bZbdKra8S3GU1cuw2SMuP2JkdHWV+6B5ymjrJTZHwzxvRQOQSDRg
Z23ELDmU7ndZkkSd6N9AOvE5g6VvRFduvLS/hhJxZ8YsK8RbV+JeX98nse3TcBYEDl/uKGXzoGQ8
OcXSrbhtZPD1KuDnT9C0eulvAa8vJu4xJETu15Hf4zfHuU9+slk35X6J+Fraun23kPj5sqTfCx7C
7RoR7MmMCZHUiPcSqj8Nq3hLlctDMyuOLxqDkPPxDcNHpempOYhP2Ez0YV7+eQ7QS6aGFnm7LblZ
X5SUZQrjl8hyMMoWQg1B5CPZcRhoarU1rIaN/vS5jIoUkR1z4UMhHf9mj8QdqF+OEEu3eFMHAe8B
PbZsVXDsUpyAiUDCSMIbisKkEJ3746S1xpqISbvsMIzFAQ2BrJ8//qUVOOsAplygCaqHPvNXP0ZF
rJu6hSB5MNK0hoIXzYpUrMANSeIs9WCe81WgQ6Z9467z1bJoD9UtsQlE6kQpL4Q6jN2No08SQIcn
gFN/q4D8F0BryJUaku1zYRqBJrKRHH6rSzztXeaqhdU8gCbaKvZgNhCKuEtrbT2G+IjfDdqi/C8j
zb8H6Iv5IdSo5uOfYauXFr53zAOulqn/yVqRU71OAkd2+PlJiCu9RVKRtGUKuX5elJ+uWpfIdbOb
xWaVe4lpCjG2bCkvG6OnC4WBka+xdnIhrMgbGjmlJGtp+YdFOR2AOcy+APkwCmxIuXU0jos4aCHz
AXXJXvDGy0EpkuSo3Jdsdxh10RzZJL/K+PxSBpZSNgXw8groZL4fJ3+NqeWaK+xz64BBtBl1jDCz
wQ7Ztu3uk/+5IjXWEQqjv+Yppbv97l8PHz2I8dIqE2iikZK82n7rFUbIwA4NdrT2X5UksYyxQvDl
utrfwd1EI+NvM6LfbYM2/mh6BottkC6s4igJcayaYkqn3zjfpzBaI9rpkGp7J/WPaawY/kIQwUTd
WHkZQHgeGWM3oya48MqsOKIgPanUUojwKhj0lfL0Eplpb8ikYTZ+GbLmqjdQMtUemF9D3cuVwLCX
gd3pAL3CY3EdUKj8EbscnqI4r0lFUsYqPGB5DNyYStOShzjbk9llbNc5YyfJ4OgXtia9MsrhQT/k
LSi8TLiLNNY/oT3iB5MTsMhRxMjtKf0eYl6tH3OVYTE4f8V8zgNKQbTex79bQbwtqxjKoal7WVMg
PA5YyLQaYUGUpXBg7dlT3NwX3wcuamluSI5VkxDa9jHjYxRztAXonyFHQ+2cutHKcV9ofg19e+CP
NCjSbZYjsVFmqXOQ+fjVjoywifUfjBW7cdSbCjers+XcCkFd3x/Ur7uJlJgbCrPC7KN7ooZvvLlI
gSyX6Wibckr+cCk79KzNmGr1++JdtFSeHawOeIuRv/DjzOK0FWQjzn4VHcax1BWC1VToMvgwdKKF
qyAKZS8AgWk3QUcWJ16hOT2+diPNDFRfYOCuYB+jUlnepcCixfPnqWHY/eCVMR/OTlbmu5wslMex
91DedZ1MicVefbo6XZuyNHDdN1aC8RhnO8BCR+rmsbsTOj5z+LA3M+qjRKkuk+SjqJiUJJQ4ova0
W7mDx9ICxssdclSQsPz2NV2lZalqlTmvvZCLB50+XCRHlMHnQFjESDHyJrHOA2jg+OLTRlMxTGDh
0BqjPcJnKFfc7QeVxMKNIsl40yg08WjDZ11cBICZJYd9rxWaXZC4huISDWXm3qU5RpY+TDoTvFRZ
tb/7it2iR/UtiWV7fzQwJUfs1KGZ/qhgVkSKcMw8q56KE8MZVEmdkkmE7SuiFpG/rC/SLYEpIDav
AGNLf1rpjd6SiOMtkwdawQlXOZ4VTEAS2Fny9MpkGwKseJ1kfDlVv+Obj7EcSjHBxUocStsdGwqu
VsauJBl02/T6I+Coo/Qg0s74B6wtS1zSdDjmHByp1VQchti4XR1/OgwRE2WIDyLFlCqfYU2QCg/F
rLdeAJdSIfOpLKftsF1ei90BTzBrAPR84aF0DmeMlnAuz6dQ1Kdhc1Tu3CMKkvOy8Tzx4IfZt6A8
rcsHehfXboPmHibbNCtQWx9DEeKr2Qrv5LxULtnaKYQxqaQX+ZFA8ZlNZHDJ1jCLyU1M6dnM3iuv
pXYjQ+tkRXUawM3Ho+GLhb7lbmBuvaSmupQ/4rD8EpV7JVaMWNzaw+FKNecaRdG6FhSKlI44iyxg
RkBdkdM/vy2L5ifud6lqjkCVfQOWb0X+S3tBjR++3z1RkEQBkm8H4nSFNS1CR1Z90TjMdkWXD8Xt
7ZBkNtwoDw6T6icvHde6vB3GneCZ+8JxjIR4dPpU8OE7FMK9G8bKSoWClDldv7vk+iAul+tdD7+b
piCcPwJDdmvDhgtQuQ2u+Q7V+oA3Ur/5PWANRy9rONc53JuXKy/J1dwnAi1YBP5CuY7hzS6GsBuw
MpxcltPTbjYjVd3Znn4YJhBiQvU2R6bSOLbhTdTE6D2FxPpeF3J7BFeUIOUpkX9CSCN4fTpNkYTO
13DbjzeTz6SrHXEWaqRNPUWukbzL0yygb8NXiXmPaHWvc1alWQ2sbnrDr4C5iN5TzO0fDG7Lvu7W
s1aAmHGbU4OX/SBBV6sgawChRdMo+SwWFPbGyDyu5b0W9afTsGvZlK27r1YlXThyJYOFbpAIq8vk
UVXcVxbRuCYxfJOfu9HNZwA2qIjkFlKNeCLUr8TFM1kyOdRLwZhSrjEDfGdK7UGCBbTwmJ+lOxMA
72wla9m9V/nOuA6LcjHBXqsTDjqVNztCes9l1fu5leM2VKXSqbfuIcgu5TDpbTUQnMUlfocLb/fX
EtsKkgJToRykWzA8cISdG1EN9WcfbLi2VqkHb7uhwjDw+Plr+Wjl/VehnZcig+lImcN97/yJ2Jiz
kqHUSI1cETwPeQeNwh7BEeV6xfttbD0QKZGxE+Z8gH5pAYFYpirLY8ZQy8AVIpxIfoOCsJrcLgNv
7OyfAtBWvke3Gc+S4KP7FXPIwD0nFkMKXcYH6GRkseCBzsEZKGMZcjzMQCuB7CXg4ApnzgFvN8t2
lYQV2z/xJuUSQc2IR5ukAaXJK5AhlIZAi2e5ldf9NeNA5qhKB2EVhIy6nrZYunadi+LqrRsODNEO
pPCrxbO7WiC8fiRX4FWkaXCobpaxVbuw/WMCGZYtqFRXdhxvmJt1OBKQNZQVVgg8PnDVCC322ZqJ
GZsBNyeiwCM13ExMMxC5eIVO1b7Csrdbs2MQmWuUQQiHEL1zioB6Qn8okSAMoovODojtPDYGF8oM
E9t2yUXVnbKqCHhHETOywH5j2y7ncEZL8FCabJl/UNRkFEK+N+OxWPvHolp6zmTZFmAFavn174vG
Y9H5Z2LR4CIYIk4fL6SRmZctiErswrNglOsMdFftmDWFZ/sMtHDVJX6KXWaQUer1PKSpMe6pZB+b
ZG1qbCHLJAcw2o42+ljatBiD56yxPpqnkE5gG+MXkalOEQdLrwxvGsRrE49VkGBxRwXJBQl6VvJ0
Ntn3xHhvKOqpOS6q6QuRUb+izA5KMvQqZcWWrM5fE+FOa9dky+rtq5ZGRQd4+V1PHd6ND6XIIrsL
SIx5bXD6CZF3e+KMv8tkJoF5IY/3sjQ4FZHmR4yw8O97bTkreyd/td0ifgLqeUzwgkvlPKWg8aJS
PYM6ORxiVqupYSfpQYUlbzXhh2OfbG+nnUBkqD/ox6iw1Xmr9OFK8e9yemmhR2lFdOEpx4czXoRy
rnmlTlxtVF4YXgbWktqY8Q9HT62RIfP78zT5F0pd5b211vH+MKkP8/HzO+YqmxoafLuzw8McWeb1
dD7is3vYyQhKOnXXYCmWIlS+qdNSUvQixUD7Ale5C0nfR0+NHIDSjedvMgqpoQLL0La2MxuuM8FY
qq9jAaBQo3bCUA3by8w5+b31vLlLCEvC5w57JkErS52q8+/QLZqPgI9kfMY/YvZ/2+ffODyoHF3w
IkmmByIG5ahzYaboK5QDhZjQN+a01edS7hT0mBDSN9wupgOW9iIhuSC+Ig58ZwC/6nNUJHqVjeTt
v2Mck7vV8rugOhF6HEJG20wVdOIBV7NkvV0qxthgjLESNmQqz9CCqjhyRPJtiEbponxh6oTLddqS
CVGK9xrpGJWA0DD9knsTgnEWIdbpksZAUhlcdCBtM9KiTB+g6LYpmhNvq2MiWgPafuoW1w/RiaaI
Lf8tp5/+45XvqamKmH2NOjqtDOtWJb5EYjzDSJYxtyAclxac8afVBkIUsdHODmXX6G8/8k/W20eX
iUTQOCX7d1Qj9hZktn+IHgmk3eUNWSeZCuc/kVjnGM3+9Y8tYQQJBWuFu496bcENmbo8Fi4ADaBz
9kESgszaDQw0dxHITmEE47iGoFdYKFw8cT+kJSrfI+zioQgp7HO3uzd8TIF63Oaw2kct6xoduQV8
xcgNNqVisyuTJREavd/lLbQMkSXwJrLgn0X+vpAKh2R/yg1g+p0QTFVsrTCIm00RUTZPKqzK0Zeg
YquCej75Gv61yfawjPKXWU/bpJrudRrz1GbpflLsG3iuAAJzZ5BZ6gqMj1EjTyYqm+pVf3weUtAu
MzrNdZGbOcuLBF7WT7xOgoG9JaKX1t7/PuKs0eKjQA+2aB3vgmpAHWr/SSdZ/tGE8hD1VnK3iuni
xhuIeGyw0A+Yl6SRhCmRpJx3i9ULD/VpKKhcZwWUgOt0Bhrl4mBizaKMBZ4H3fS66sbUEAH0Er/9
5fmcfZJEarHeC7QZ7ueq41ZYMoD2P5JSyZEptdBaUxii6LNMzw5DDTMqV5MoulxtSdP9Wdd0bf7R
WzkM/OzwU/r1sIDljyjKgUD8Icay2qRQ6m34U08EqDVMgB4AuaHgpaVWf3V92aAYCrHmcw/jvN2g
gFzUk6bjPXNluZteN9MqsHtCym2RuKG5NvJgaZLoOwASvWr8lJu/cwHFSkFH1oAdawFhgI1Or+HM
cTpmeUlimbFy5h47SJySPMBkYTkZY7MVqz/AtnR68AKOEVKUo3V8/UKEp4Bo9Wo1OKK7aDsM0OS9
2QcEDkOwW/dJvpFmCr93dsRlNzsJcTC96Xj5PmIJxtK9SQSOrNuT1x/UwgthV4ZdNRX/WiwVeDYb
yovsfmRuyWcdYTu25sqpj2XBACigAfEV5AfW6diBjWjAkj1vhbKVich1p/Vsuslqsm60yPw+sVrG
PLRbdgfo8p3xVcEUn79YAHFMcP+6QJ/Lld491/I7OnMz0m70p2rUOoEYlp/W7e0C8YsqL2CpLb+C
TKvYao9RP5VjsTB/b2YY5wZYzaWmsieVR+NRo3L/VgSZFrj20Zzgy76POFFujQfKIOYp3ieShDX9
Q3H4KTKmMUpHCKY1EAPIO+g3Pq2oAOdmuBzyaZUdR+8D3UKBI0nA+ibPAC7bEr357bCzfrU5U27y
f0sG5NSan7cwLooAZU3FqhqqzpIQtzrdgCMsNvFePFf8lVQ93zdRz4t8+gVmqjGSMe6nOdmQ5MBt
HYDaIFx5hyEPmy0tVCXMZZPHcp5xVzMtP68p2umyKqhWOjKXC8J/7K5qoMQbg1bDojqgzlUE3eaX
96vwOhQEq28y7iV7auxwjvKVsL5TJyAji/Vm0ZkZPuWKSc8ONPulDL+Xngq7kRgb5MYM3mSK0ua2
86p6r+NAIPd9oItZWN/c0kK7ld7vfe9Burwwny5GEryPpXcxa1RuYridXCNCJEQxKTkUhaW3lIyG
vaQwTu1Z3e3bb1QLWCnR17PxQwtXfQgjJ6apK4X8TAAypbZ4ztItBgI8Sz9/ocnBLWJoR7WuN1BR
czqtaX7KlW3/sWYz9JigaNSXm9VfdMLsGqFhmKwd0HJGGOF2HaVJgPxiVA0ScRtZ6vwcW3fKu5rg
nEgqWH7W70ayfTtjY3YsRCXj5jaiUjPS3cqiyFQLkgg3tXDsDRME9/aj8S+Ye2TH3ow4i/VYN2Cl
7O2ZIxfXcBTaMNrhii/7rXiXsrYl1aJgNA4qYPl4VZCNUZdXlkokO5E81zh2YttRMkinOaXiaMIG
S6i04jhKVMeghZejkQz1bqnXhVo5z2Ew0X5eeJ06ciQx3DW2gq3H3wpzdpAFmPPBm1EghmYf/7IM
TQiG//HUkGJg0ZlF8qCp7kjmlpLQ1mWMpO2tPQRZovl5Hm0PhQvxoRxKT3ZzaGPpihfyZJzplsim
HBsFoeM0/dii5ySmb+f46Zn/+6ZpNK/KOP3o+K7hKtkHe8O4Fq+zPaMDZtRuKUKruvn9cllGqUtI
AHcdr9LnhwdixbHAjGiN8tDiCxxVdpHga+IqTM2ysylVE1sO+AyELCJDlKF161eDZ2MYkQhpyP3y
+lEr6vqIcYzGwc/6v2qHM/1hYpc+EpChdYilG7/F96I6Sq5MxIGH4fog3iKSg8/0QQOW6sQlTgBP
JTRrxe/7oxzGwPtHxWr4t1bhA7bIcrjo0QTeCj2CGnhLAjzyqLN3KGq9Y1uyKw9uiQLupOOYuf0j
qGi3j7L5bAoCVKscFUudRlnJ2P2Q5L8fkk5LJc6pFSrzysvJmokCA4RSanAzT/33g0aEh/u1fYAp
enU2OBB7gVvOp7KWJ7BB7skvg7CC7S6YMggvlMdTcwZ48uEvvv53e5PagUOdPVqpu/zTLyrAIzR1
sctq/CLQxJ4Ymr/j/Em1S8ocSdB+kdDnNSS2UAvqpXc6gcI4Cf1t+CkOag7lnAonLhshYbUavnYP
4knHGZ8ewHEIbM47pCfKhCh3Kz6YwyySO8hgoRvrmKLw5VclynFiCOO7wDrVOwCEdiG4ETvuc/00
4ITQ3XRuEArksdLxjEtxA7w3IArfPMPGTRMU/lxu8H1BKdNYqzHChj9cmPNelQlDj4XT77OUm+5m
I7bIjw/OurQ7A19JqcO1ogp2tD2tTtaPLqahPiWMcH9hWnpJX+4VS3qzYsPCsABM621P5Tl5WEcb
WEsqeKiBCzVlhqmWBz/srageCz0c0XznBoj73bZ86aM1FgjeGe6dDvAv9blLyqEHh0XxxYjpahU4
2hzhB1AifHz+LZG7TxfHoePQe43YCGiVnaVnozvF/hIyqobxvZ88yRhi3LfMqPfd+v+X28hfMUTS
n3j9O8bddB3HJEvziJPUD4RnE6kKuKEM7S1TxgljHs/l+xwNCWte1EFCJSEJXaXH9Jud8bZPcgMR
9sc8J6RyJiBAFcN4UEVMqcnp4fhpPs+wNtxqMdtPt/ukYVQCMbfwYlwwfrbq5QMfmn5Zez3ePSST
izOUSDOFirmy6euiKtm+ywQIM5h66jTa7N8l2y8dgw5rRII5fHJQWOVZY8HRTVMi3EyyUI9mPg+l
TzCSIebrhoc62/15Sy5Wx265zhSbrYz/98kgiNMzYX4sVKqsP5AY+tfOswgmGyte0qOktTGGGOrG
Qb1W1W53RF2Gs+XU67MfnumXF2AUr7xdRpe1EvReqpMNpMsZBquS7jJ4TWeb8Gcq8I5bF+TfyyCW
KPPlJeFOhI/sss657jEVok/RbNjq283z1RUbE8O2NGY16gXh7QEqAHzAFNIwi4tB7Mm8lOrtLBjj
IzKcKQOEG4sRig0OfnHF9DlS58uH72+Z1SiUzAWB2a+UNZAyuMEuFD3lPOFLblAND1onraSdjLyO
qZcTuw+QqgHXG5KUZ2JV3KaVoENzreRuJFW0kbRGoTu6We68OIctCNeplzFskrJi6GabpxaJLmBT
6tuF4wH0cJNVSzk3ztfLs+DRxcWZEELO6N+ytlL0tX04x2XELHLx+BT3v3IWss8SIIlQ2kvaR3kn
n0mCt4cpSItTOg9oh5XE7W0Ou+IBo6UiI2Ytkf2dDFIpRjUbOgR2HtcebKaMlvHhE1Cd2CPiyJ82
FOfgb2IZwCLAGeajpCSpql73mZhYe7z/wvRikX8Xc0Crqgw67DZG3DNqIeBZFunAyI6LSdFUhi7a
t/nJMe43LJ7+D7YJEW6LZ7jDWFM2w0Su4RzUEdakD3JKiatqtnjiH5efwGJgu88MTAEXlKfXVqrN
q5GybPUuFbRhK+z5ugQmlCzr88KiqjNO00wj4AW3etAU6dVBy/+GMMIei0syN3KY7WMbbuQnUJKq
XdbeKrnb9UPxYOYyUKmzVMSsY1DkYbQOH9I1ocxNmgJURkmtLtcRPUp5lDwcVh58dH2kBp2Y7ANI
mEoTAA0qx3Y/KUQ5biubwRYdFDdvEvQmJS9uRiMeCnk2NWlHajVknRBJrA+V32eOaqtGAyszd9j9
Wk342ihul3ud/Buevqbw2/Yuc1NWwT5v4mZoRMmLGOUal5cQbcqPWmeGzsNtfhGKj4ZUymoqgaba
9JkH9oaERdsLcvgsnZWGqmc2SeKVxstgVC6l07WsBDZvinLUye2Um2tbGh1kzO0LpI6SDWwQMkUc
fmPgjhqoj/dGZWYetfNTjXJJNkEY+Kn2vKO/Sq5zaU8C3Uw6ksbSP270Bqb0crmnT8LYh1dFGud0
mdzFwwou22xnYQ3zaiyLOVk4/uZIoCjdQNLqy0YP1918E9E1/pBThFxEWQcOqZOpQLxMbuI8cgS4
jcoAhNXK/2TpGrg7j13AXMZ2A0RqpN8cfkaZ5cnsx37Oi7gQegYnUwve+4V9h+YrAxrF5EF/kSrQ
MLQxlZtZ+yV5AsKIw/n9F8yNjfQR40vGewMouNR1JauTGT+e6YmNGDUeCVakpeBjaV5tDeIgmuaz
jj2U+81b4u2CeK+BXfLoecSb98fHjmi2fHqk13+A0sCKYfOrePA0N/Ujaeo4MXdi5AnrFHQjdc+A
EjEvNRspE17jsIMnTREw6G0nnFddTjZgKhbKbQRjxgdCu/PuQz8xZixFtiAxhANzjNhbQ2tGc3o5
B/JiIMl0CQZ1Oj4s++pEzBHtWMjs1wG+0qlEhTlh+ZFzDRj1CM/pNq6WSh8/BJDCXtLWva/SwSQG
rU6LxYf08+rl4HEn8mfxZtaAPCDe6c3BppW7MHwWQL5WMeLQ95YaqtafZY2y/MZaPnc1QBG5YyDy
YUUehUM8c91HUGPUe9ppdZYoAnXMFDM5OsEyds7I6zB3okLPfwPgNCARqOvIf/jB9mK+OrytEHB/
ycVE5vTwqzhwFYOLr04cKKA3i2t89poLs+AGevIhJPuzRieia6sr9619sZEgTCGo85RkwS8XCGxF
8nncbOSgHOabzAwTnyar+TaLRmt9ez9nfczKJri6sxgKfo5YtUTeH48cO0UYB60nR8U3/4HFrkjL
txUXRTVt3E3AHTmOHm33ebk9/n5B0m/n28Q/bCxtweoYGiA+hJ69KgoAGLHNWyqlDgCYrV7OR51d
MYhBUNghSFN1T1l1KglECkU8yEZvcqgkroyeSjcV0fYNqNVxgtPUjGVe9OK4Q9zjfzOWrz5SgQsD
mKwK0Ex+JCjPWTZIk4gFTryvUJJ/8L2wa2A/Dc0gN5HVT8Ku9lzB7vf75EXMart1lx3m7DeKlt/L
389SEbBfdVBTejfUDzXdIU5zB+QnhFXW6bAPdHraEf5LF/fmTxoPwHRmXKi+EXC+Fy0uQT38jd/L
4M8BBdI4ErAt4OAdYVNeaXleMajG40rF9va/KGQrQlTt8NKmcSaUr2JCnAR2GhBI6RNo48rOlK7O
Eu9+78hPcDxYQPa1H401cmE2z2/anMG+p9FTRCr5HfwKfhQCwBd+eg/WAg1YZBIF4ahbb94iLb1M
MihhK0BjfsfoPjcFEinF0fgpcKgHK+nZZkjJc+ZBZuh7EOzI20vEx23eWd3EcoAiAUxshdNipNPq
cKNE3k1rsB9W7q5X8Kpes5eLsZ6hThjWz/bE4ApevnF3l1cO7fZHhNunc3lrqZct7PSOUqeJHaNe
dfWDWFYx8igcZeTv92oVGvmBVyNemK/6OgdgyyC8EFbsZDUFMXt7mNmEPf4wxDZzgMQWk9wn1SPm
TU1pvfRCuuImEJRqcrRKU0HlYm2JiTnGWG8pcc+QAOqOtg2HPxfpdAejiFMS4h3RoUjAX1lSuqZe
eUr7uiL1LR1bqnJ6TokS7CK2TEEu91WeDhAvm4KnoypkkBGuXmefc8TLstUk/hbvICe8dmConkvE
YuVAMrtgzKi3ZwsopebUsifD7EMt3YAU1JKrT0DSt1XT4sHfhgyq/6qCVRrk1D97psYVVYg7Hf45
ptM1NrNBYmDe1KRFQ3cgVGavmxLP9PzbeSFPicWcfvawsm4+u5ODAWGoNsDAhZX9e1xq9T4MTU13
UthD574zW0zkavKmjD5iRvnjpDvpsJ/dLSGYnRrT4nNu6PhvRMmHknK7dN0FZnqmchYeaObm2JeL
HybyudMpnTI1MpuCEiYPaHOfmvQaIJjXdF8llW0LgJkhA+bqafCgyxLSqcFPpNSeZOoevbuyOpco
HB1L5zHnveA8tKScKIJCiRS87+hCrlOP1ZI4xl+dn8mdvFWNzynOOYrw0xfAzRLzkbA+NYIhMQS6
3UUtwNFFJhTcdzAqJ0HTXDCv/wJqxoBvBNQ6xJaAM25T/GaYUbp/uhvyl2O/Bt6FMu9+23oqODpj
04+BiSkjRiDaTLgMGU0yfpr+gkdOfHaJK8jwC+W0vl03JK4UC2t5xHEITjx58gvcc1uiPkGfKlPL
6GX8EL1ZgTvhtuUTqiJUhnsy5D/1YBZryBFZVCb8nQpBjRio0eijWBM9cc1R4VyEaREfXigZZlTA
NViqpyFs+Hay7nRtUMRHzZmd3yto8xIiTSpTtbIZlZslx8xhSz9uUYz76KeRfMRUcbr8nqHqnON6
taV2tSmjU/9NfUyIGRBWnXceerPU/3ok9TG2Z18yaDoH1+tOpKPdadgNSA0Gqz3nUIfKb73wVeqB
+4GNOpsCN0Zhx90g0gximQWnGBLgegXRyRH+SOop5HPmc9rcEPjcYgfWbJI8wR3Hagskr8Jbc1Cr
DcTGpsTdLOeYlo15YRKVm6PlG7ypZxX59ItB7LylS6qk+vDVJRM4ajuTdiOb6SIIJAFGwGYfwmXE
cX0R/2dbriUXwP5AzLt5lRNqDiv7UubL9KndeIH3TCBqgmeaOjP0IHtohy9yccgijNJvj5K6xBrZ
ilvRreFYvUL4svJw2FPzETGs2ebxvNQSKgG5edQoMV1/QsHiOPaJY3x+hhlTrNJGVPOqiOtSOsKq
ciocc1buLdnh/jfkwBWavjrPTqeQF0vp9mQu6no6XRI45nAd1R0EUOISas25ScFK99qJ9ZpQmGbV
2tLXRgQAcJyxCycRdb6xgZ0gV+6DNBDwIklwKQE5iblglvgWkkg0r/tAuSBm6F9NN92GT/VD0/oa
uHSr0hU6bWO9HFy8MoSnIGs6JrFVAtRuwsK1G2hBQBz69t5vGm7ni6ZTFqshSacPFFhShimxRQTx
x4j+NLIYtDb6pqFsYKWwoB0P11bl/ubfLEuughUVCKjPcJsUcoa8e0X/wA03CmsxD2/Lata9UWKS
jb2TEZUjZSR6dIuKDt0e+k/MOjudqrDOXCwlzl3shHCqNmZSS0Vo2zDDUT1VXqAP+Af+avjulkdQ
Dw0wTnVT8MJdtBxfQ1hHS1emCoeBqCLuGuTfE2Ud1Jav6YIdBZHobUFl39q80naye9V0ikc+b5SB
SEHmMmy5G7knQWZYsmXHqWyzooUHBguhB89nJEXlux0cWpY75pfAGxlhiMTePCF296LSlOzo8mOy
ZLFgTwtf5VeJ8z2sh9WrR30KR+XjulDMCFEFKszODBCdJeuaeysiuJ/qbni1VqZ9XXdJ5NUYlUE6
SLY02/+zr/iXqINzRLbjSVFBJCUWJK0a7XutsGqaYTe3ShAGdkZxaMjQ/zyAutUXQgoQkAe910Ep
hC6KZ/zekGdxf5n/LJlRJs0QkBicURBlKq7/JygUcKlR3Z6batG3UUrwnaXPVMtR5e+GZqNsyU4H
+WAfItWI3CUbFPwztXeGo5NniJT6k+oVtWyaFZeyKYd++P/1bmB6Ndd8SbCnR265OpVn96H7gGwA
QgOFy583ip63jCI7lZJO/7VVavrntLdjVy/gKfmAaIh8j0NwbZgzvV3ErKshPOo1WZjh9QYLdU2D
VmS49YyCvPF2KLuaqPub+GqESUODKRXfKQ7u+zmVZeLKJ5Glz0GwfUdQkY06dU31E3FCCsaSczeF
0VaI/X4KF7FpxlNaGJ+RiUeE2AmxFiqZ6cmN6wSuYTrRGrB+DRtZcM8EzcdPUl65f5nWtc9edKeY
xtko1Iba6tMGFA2E+2ihiopB7143xQQNVi1nvMc6jhQKoyZpGVRD+1srydHp+HAJz/nBYkpjlZ/H
QHnmudGIQrl+1y1O1peFBNW47Hthbhbwfeytncdvwvoecu8U0wKWv42yBZsXBGvHaLQN25i51xi6
UtOYXl0TDgOEox0vm1OKBWbLxYqbeOnkxnCIw8ad3N7hj7OPPJs0bUz0OyDy4O+2ClVB6TKXHPuK
KQuCWq2V+cTrTycjmQPdP66LAy3B/tmM9jrZqne2rSysxcjGee8z6JRX2QCLLMEX3bO8lKQM+LOa
RuZxsbkJV5aMMbZm8FxCZHjF9lJDkOphMoQhp9sjTtcqbcwW5UNu2/q7DtJyM4mJn6xclqwKXwC1
QY3AzcQWMGbWQldDVt+aBH8DQ+8d/ES7GWHlMkezUCZrMx3SwNC5MS5grEbmZ9CGKOXrN+jyg445
wt4+JKPi9trF0I1ffQ+s8FgOBtDHSFx+talvOc2fq0dttn4zhiLna0e3dRbOe6udZ2RQ7VkOt0wN
nJq+0sYP4uusWK+JvTExuUSSuTZDm3d3q18L1LyKcshmdifhqlwzID+6d6/SYhV+JK1snql0dLbJ
lPl3BwAp6fHugbMrAVhOvdZQWHwvPTyP2Lbbhm+ENOgXd/TllB9xV5/1cQ9TQ4k5F/bmP0Slkhw+
9UFqN2MdQaRSKc81TevK/dCpxG+HXhN74f+wsVA4unpR4rz7jvyn+r9vmcuVza6h0xqyAqMESHRJ
P++ZSKku0V0f9BTCVt1Y4cF2bYHbvcaov/6z2vYCwks8cwnkvZmWNrFU7whkTzun5Z8Rdr+72MGL
CCbRQxmsPt7mZZIHijcwPiQHjc/pYJIrajhyzXgPnzmeTXFYDR2C+iv3XdJ5OvGzciqNrQ0dxJMj
mNq4Slu4NINhCxUGvi6zwUsyDimjku2xGTPyIgco3DR7oZMo8utOcYTb2ONmcdc1n6cKtaQGD8x6
ay6gkURTFYDDPl0ficBVwAed2oV5T8cXgGnL+VcLa5qxLIgaFlTidI90Ed/6m7DBPvEKd+PeSFTW
f8syRIUGi57PJOVCvzMJQ8nciJJgnWcHQzx52PqDKUPu5Axwulupb5pl3PndNMEojFhy+3z6V3Ej
hgKcs1QTKtKHLPSZJMVfqP+Td0m9m/0KgaLDcgRy6CAMCB/OCixUa7kqnj+p01vYhhSxNLHJEpKU
7UvgP5il16T07KB2j1c3g/60InPEJxMnfvcu9eNoS+2IYCKuKBD7fAqi/F8lVYc1Maj4KDAx/7pO
Z6XnmdyPDPm3DM/PQ6gIfeUOQV/2s7ZCgXiCp1MiOhKOKja3YnR23P2yoJeils/ebjnzbt7yrTEY
/0xQyP+PiHy6rGh3YK3LpLXR29/TVkLri7w9Jj26NLylYsF8jPlL0hluyBtVWa4ZcBdfZsqTNTHj
W1i1cm4GtbxTiXXA5POx1z6vsufD5ODi1Rk/hXAICOnUCeLnfWASOxLyHIaD9pCilva4U6FRLv5k
LDE38uI2OfAxfTd+3itzGZ+SMaKLcH8eLqy9ikCL9NhZ4wMsOWqOQF+C9o4GWXwaqTXu/2OulNV8
UbfATWGWbdmcebeHBMJdoGoyuGXzA5hxbWuf/ZCz6y8sDszEarUtNegK3hO/qH5+qC5GMYH0eXZu
ms4uOUyqz5ADh5Izv31VAwkH/PsesSBNt9OWA44pOJ8CFaUFDTcL/Ac70Kv7TYNCHfW/nvtRa7Ri
2VXqs0vn7qlvIXy5WDtHyOwMbcchSkHTRYVg8MmUjISpnm6Ru6dpNjrRnTtwkIZuw4RlvvBaadT/
zTQkmLrEp4751XQoGGXikmlI1Y4Un+5zWstjtCUq6xCx+Q1nJYdPJ7k4oJie+LKHnYKcC2t3436e
li2bLXzL7XdBqfyQoiAXTs04gnUTdWOh8t8DEMK+ue7Ow1eJIMAVCAbrY2K7Wc+YeAm4ypJ3kidQ
GbfKaJ1t9KL2LlUVGSH01ubzkmuIMOdCW1bzZia6vb08n+CTIRUIyDqhYqbd25R4igkQS6v/BalS
DJCfLGrjlB90r8DnP/PHrmLOQG+paiJ/hj2GLreShs96eiOB2o6nzBGD9KW8rGu9qB4WEE0zExb1
LWnkYFpwzEDFTVsQLNDFfB7LOwNntq7VzsXvtcBIQ9Aw5E/lv6i111uf/+JZFQtz4k3Y/jABfSBi
7phm8VZDeD9myL59mEGn4P1q+nN8ojz8oVr0Fha4mUMQRnjLlqaiXGexzGHI2dftssB+wsnOyg0T
15BK6hOOA5NjXtDRbwp/jzzsmjCQPIUOzhOauwL5SZBoN7Lz5ATLsgYHoovWgr5G0k1+CWUIbElE
HsAjSpb5iirGOITwGgNhgb1uHo9ZoxMYEW+yw+plCoyYlPIVMWc3AAjm7cCBgwh0dy5ACkyckHhM
dMKC6sSCE8Cq0GOWVO8EFXnVk1b8IxosAa88mbv4cMRp3Vm4DMNiS3OgODJbkQXlvfHxXxN11xBM
z/QKwc4P9+67JI8lf7QKevvHJeO70z47U/J8j+wt51U6v7r4yLBblPUBz40qoSb1JPvQHdLB63us
bSfsQVHRHGv7kanWGW7PfDqJVjq7yv4m0XfGGP6Mb5kHaPN3EjMvpwKjANaMa20mdnayn8obryLo
z1it/OICNt7MIcbIUHrP8kBLiMrYTeQzxQ0xe7vfUysxojpUsMH5uf/HJ+oaXGV19/EY/7Lg0+Ir
AnlMTDNqAWAKFL3VZIRGzhhfs91Ptwwsdtdkerv00UbtK1WRf3VlQgK93OHHijaoGHiFbBYIgWd3
dhjBtiqyPFvawbxSuc8qpCdXB8nDXpsHu5AeGz1o4Jb7/FivEVpx1u5WxfO716Sg+tNseA6Zi4P8
sOJG3P8HNNc56XoOTs+URVJ6hA8TWPV/K/f30J8e6TrB2UuArwKGyO4yap37EsQb+ys4T79javvF
8GqyytV6tMTzc3HLCJFLqH7aXum9EdtLvRN8ooQkTP7tC0WjWHcrxye39E8lM5J+LDSNJwqjiN/W
moqggPgrPbLS+Aiz1iBETyr8+aZ4hWR2kGCWlW2HFNwNu+ohfYP2CLJuKekyiICqY5KyzdYjstsB
dEpsEeGeZ0G8L6/d2CewG8qH4Fd2y0cIvO9oHYc/5oEceH2TFN4+hIxg/dnaofpbFfMvKTkd/EoK
UydpyYnmjQ+FJdIx4wrJGpiHzRTfU4febn5O01N5V4prhfpi1JXlGc6mMZCjXEWWJRC1vtdMweJN
91HKhWkENPoflRnmXluApOwQbkU98USwrRjny7c17LO9ib/FGYY4vNYk3wIFb9RgmgHbOyAw4xOb
WfBK4g60e74XL8Nfz321bbFJWCjslLnGth850K9rfGYtEW7PgbsAd8igQiKofRDljEGLjiGsR5xn
RvlGGGax3Dj0AR9fxn1Lb27ucYYwWjBBCxBlYBPHSHVET8olglNodPQl8KZBw3rs6JGWxHh8wqVC
h5Q0VkETe8uEq75S5tDKJwXWwI8Jafv04oXxs5LePanyyRI/V7j8Q9Rr+g6ksJclC4IHZAyi1x1h
wQi2atDiD6ojvsI72SJthPyTIED6R443WJoRH31rT/LxjMO4uVX2EZOETMjcoSuIj6hVNVy+xiN/
TRHuhgZtWwmDsAO7WXZE61FEg9VxjTfPTeCfvBbJe1xL4cjZWP2occaYPrJ6BhvOFtnAy4w+QU65
w7FUCa5mI8gOBA1jMAo3RJZdsGavJBHA9KL0de/VTJgxcpIzPI+iBSxBWJEAqyrmqtjhUFGFbRmr
zKNU7YIoHLLXY24sTTmC9qtw2dQf7V7lQWevZN9VcPNpteptY4HbujPBNDbB6raTiTdkWYW+VyjF
HytR25sbBb2pXJpMn1Z+NX2mhUZLbjvlBULUBGoaa3c4oEc5LFHddgX2uYVxTwt9i9bItifQxnuJ
N+vCb26cWCx5g+AEWJRzpaZHyrfDdrc3hEW42Wfa9I60w0eWk+7pFFqvAE18inVw9Nslv8efi9u7
WfJ8K2OBi6u141/oDrdxRjCnsIwfxU7oPlYRt+1Fh2En7EhjfCrIJdCDW1RQtzcFwnC3hvMZMJ2k
f2mhTVPi+6LeESoub2NC6SDXdaTbO4kKAfoPLR11r/L7LJpbO6+GR3AsjWH1gaRMtWxO983kv7P9
s6b+xVSUSC0tpKELvsG8JFlw772NcXDDoIeOM44NudmTAu8wvUrLMhCXjxmlvf+9u+BuIfKB74w/
TPfIyow/BXLwsvxdRdjz9HgmhrNPr3x78Y4lp+2n7A4jXr874zcDeDTN8zH0v8avApVVQ7CniwGH
v0TypHXlYcOHYdb4hVavnVNTyn096a4pVwp/6pSVxCzShDinFhku1OCayFQWjJqN19pvn9uT/Z07
g+mVz8/BUxaCo84G1XclM2MSXRJ/ohSQO5CB0EjkOXxBSUpUgdaFTTWC+QCvxgoQPDq/n52OAE+q
Y2QM+Z5hy250IW1OqlFL4bHL60DZcmilc5P/5gqdkQHdOXtQ4k4jfJPGKbusQLRcLIQY2AhiroRa
c0AYxzeH3+2W8mdgDUS/MWAtNuVk2uYXksh7lO5J0pDXwYQnwKb48tEJ87rhhBdkHAnUK3wsyqgj
9iyeMRQqx8td5d5+JvuqcWEHMrVUIV8Wa1UxLliNGDf4BHZTFhJu0yYdGAt7730PFvvXxe1W+Wom
U9hO90gMUBu2uvMKye792TyZGYw8o0cVPZGBusATCStrM135M2Ciwu0X1E/9JQ2NGwZh14h03+Ux
tjxcb2IKpi2n5KgWPjsb+nh4hPTzhBlQTpgqTjnX4YtxKcOD4CmC1hF0MXG5dczFSGvMiVZfjZ8u
FZgnApZE8nG86x8YOSWwqfRAIP/J3hV/KM2JbMluAeKNOvCwGT7w3pelm5G7CfljEWGM0owXSChE
TR2kpKSymzDRRrRebxTwdT7zB8rgyfBauSDKkHWUNDt0rNfNxFqw/S+bhalJ4clTz3Ln5G4Z89yn
uzZ2Uhc3YvOEvm82eDKFflCf73Xf34vRaVZhI6H94SqN9KSydUdJKeTzKJcHOuao+wqTplhayBQg
UewU/W4IgesHJ993VkztYbloTpQvLi/NPp0rNbMrAXDX3g3dQIBCT6SPwVJf1QG5HQzP3vwsyEKp
3lV64wxISu4BpaGeZM1rpRGhGQr5El5/Kpu6Guggv/yFrgO5yG8jpUbMaJ+48lu5D43uyuXroxSn
qY0MbKj7w6Cst3PcNGYuU670Seb7/geW4wPAdiu9adPTkzfBquz95FVvacdrCEmNcBSEM2MwJB5r
4zQeq3xk45aKeAM+Qi5IOaQTBqZ6IvX6MB8CUwX4j+TpzgTVNRgOHyMobDPJ4J1CILnFCTvCANCA
9WEXqPDuNeCtoRYzL8w3JCBxgOGCSwCZdh38FSXDbbwNBB5czVUOkMp6e4y/kJlupujFUdOG5TOt
v9AqFW7pU8+WVkKG8NTdWyaj7WvF2u2BEVzbVwnw4kP+UuBiMnzIc0pGqzetSOvIMq6Egbr3VhEU
Ro5n38Q/EQPE7BmZL/slkPkkGALW2RwI9l9Xn6pBwy3vYeEoUdnRkI4Q5UgGYXgPhQ76JHKEgiwA
gnX4+RB+++IbMDbI6GE/6h8imkHTUqfaxcH6tGUDG4MVfkYbFV0LWrkDcCEDJHy4eNiHI7gnO1sF
QYSqNM7knWY31+kXgP4Rx+zappGRhO2c8WTBEvy3/VZtS2VFbaDnOUmQumbFqYf4LVkiDkMr0N6p
iypKarqO7PI4gV8c38sPlh/HmTAb6tRlCi3uRkON2p9ZI30DvznI54N+b1Vehm1P6VLqvu536LcV
PJM8ITeprK1Sp+6feBCmWD1wO6PX8XW/iE8FvW5F/48YKVT1zRq5uyjYMicdDbe2LqAHpxFYx0Kh
x2ID9MUrBgGVLsymNhTRMP+zXdv7pcrp3k4ctbFFijWnW7it4nFlNXdZQ6PW9ZLNtBNwgowHTRdQ
TeHgtiq1P/aBJgLpIFFGxa654xISk4o3fS+VcHCw3vzsZd0LxCI1yi/0JnPPCJhI6DTn3xNi1pur
Nw2QfRHYrVFYxdd/bwZgvhrCYi6CiXHiKlUCuwYPv5vnz4S6k/0/TgBmhHObpGDH2Qkuxyjwzq49
K3sdA36AJ3Hf/1OKc+Ws+TVNreFYwsuorKT0lsfH0pVKW9GQKXYhhB5ug+Z5+3Hq6VZAWTBHC51z
bBoSF+rzWuArectYbaCeQBlHHPvFwGgPvzaSncNFeu+SH+AK4qiLu4AmtqAIKT9glBcPZybH4G6B
BzRl7w475dSAMTSqZDyLVTu2FL7kNgMSaXk8nwbc3k8sQYeLL2LWIjielAh92JEk1OdKsA9mNq3x
zrtNlrQdE9Q+SEWRi1EC04WMCT97l+7B9NQMeAkVAuE/jqEnt7xt0RoDyRBoAeLpoaNsrUjugcvx
tZ9Gq5YA4y3YTJXzHC4BPlS+JDhUM5vJni3NiEz8wzSJXA4WYZYM5fkkRTcAt8KovOJN0LxZhoSB
ShOFTISOI0bwhJfOYrtxcPevZhHQ+0d/lW2vcuy8G0CYhT+7HSP3SYwItAIGmL9Ug3fz5pb59hDd
qxml/USqoNWJjDwfxZQ5xCbEsY4fCbCunUhcYAhR9LNM7lrIPlECUAvbP1BIHomuBKkb7vN5ImQY
+NlfNawt58syKUpxQ8CpG43E5mkueQmfw5bDkwyQy64y37r3BhK8MDLEFhSljQj75zaVIBS5vZLh
P9AbZr8TKaAE+CN7oHYpW1/QQdaZ3CvA/hYPi4hutjxxp4Jb7MF7QYM5dtOd0OJrzCeStTRnqfNu
rOI8X3rTgss/ZfsA35YqF0jK4Yb8h5dW0Pnm2CCVUUFp3jFUOkLTwIbqWizuI/x6mHwDK8itvwnx
xRAat3TC9+EffsoUGr77vAguPcCbwm3QjhwO35z5uxQ4KGqfkCVvag1+NoDXTDI9w+utOIxxq9Uz
yLAkMf99loQfg4fqdEVjWOJlA+EAeVmLGesWQ/GdanPodIz9WpB5n1yQrZAK4CmgKOwOuMI39ezQ
pnwA+vobZ6cQUpn615lZCHVTHD+Wt4Fegflx83qYuLoaSO/V45QJStP8cPxLLlFPwJZVBUNbEMW1
RwQLww6v01SF+C0QbeQ3qPMltOxevXww2FDXcMdwR2nLCPh54OitmZM7D+Tj3pSSU8Hz+8wiI+i/
+IeiHKoVvIMThVPYyoaZFQPVNsASnqbx+5beCxFtb24vm1ynSvUS5UF5t4mtnVzdsRZ9b/lzQfVt
UsOpMUQ7X5LKEwmjQtI2mK3FlG0obDZ8b43dGXxDMmgo9j0LhxgQ774EUa1AzeOT4aJ5OcMjpiqh
PJ0jLiPcJU79ZyYTOXe4gZ+2SayUQVBDUC/Nw3SJPqYSj62U0VjEK5+gcThqhnO3mYKK/rLyAbCC
3q++GOFQub8Vs53s1hwuORcYsKQ8/08HypPvkoC6cctk/xhglustaanpq6cAdGlvQP+vBurABXIT
T8d41HyO9Fh0F3HjvQlLG0l1eCGSpos2n3o7OY7Jo0o/6T5EXztfUEomSFyJrCk6izx0GllI+sls
lsbt2HrlwVfQxXZ5xWTpXDuZ5i642Gam+72x9ILaCGcOx9LwPai+sQPN2+MSH385tKzrOV9vS3Ym
tcrMQXE51Ybc4wRxIqv9u3fungR2OYsmXKaWWnXyXyskDowXmxz4nSEfa8Peear+xiJHa6Zv2QBs
wrjJmIqqMZq/LhuU5qKA4AtTRh74KZK+s7WGPqmq6B8PVwP3YIb+cra4HgEa5uwJcE56Kdhdb6QV
GzLFlBX8qfxU5Fq8pNzRaxaepm7dd4vLcE6daBEjZwqPKWewcXlb033HsaS135robus1QbY4CehE
aOW6uVxM4b/qznNV+sCAlJalwUAH5A2Jdr23MTb6RprIg+d2eAILKRdIWo+TdO67YeGQkTqAG5Jg
dj9YkdNvbpXDseOWxK8FRCM3RLeCxh/KMMQa40MqetBq32IApzzZ4aePnpkMnQ+7mTKDkD7oXFSY
176esUh0sexG9AaOo13XTRzRjtSnOEhYCDtUV/HELSykOtshPBzF5dCH21GBAfLDHOseUOK3Q3JU
MYCTa8eUZIG4noC8HpO6r5Iz4Bw2sk9UjDe4T/nzDXJfGGd8hRAF4J+B9pn8yxTfrqSdiOYeEHM2
77cBBcZ1iO70JXV8Ol7EFpmlxtxhysG4PveNOqWt4Lqn7ZVl4t0g+XSG+YQkbC7D6ImvyR/Lw/Hi
bOI15+VksInWuCvtmVFnqSl7rURz53vv9GNs8guFSlwchLtwLTtfn5WPdTjpqluLe/XLm7l4k/Yq
yVRT/c+3mKEcpQIVM9WL9A1unh0JkwOgeQ0SpgNm1sApCHQ6YbaSo7wEf7+tDXOnzsL5kmJWoURS
BCb2ffLbw6dWk7yvG6efZqHJ0id7v/uFRHuyOQ4PRXPYNiaLqIQW+rRxFixrCRpiGweXE/2CXs+v
jI84fhJMviEZmxWiocSkj3EZDhDIKsllEyIFzJUMPLhdHmtu/656vDd7UmiyuD23GJ1pBfoK5faU
gDRHyEOZDxoqAKc9uv3jRzHVLeUPYXGYseLkuFSjUx2D7VXbljza+11kGL74XmGRL+xYdmncE8ve
QsRTMV1nx1Hb4SC1HRTtxRpn8aL7mRY7GFQhduBI97EPnfyj0PYU3KxzAA/jSsH//ZBCm+QRU5QU
T7neLFoSnsXs0s2EGS5Xw3J+RrmxX4kWUYUfEtxqEdjhG6ivgXqxu2d6TYwHHKk6OGDXY8kqB5Y/
7Iw2hC9M5okBgb8AeT6RpcJeKKhVs/dPj7wbOcLmgjK/cNpbzd3VUPWEjfDO+UOru4f6foVlXF4u
s0pH3eRu8ALC1oGZL/G1BUjQzPhD9jap6kJWKCNMwzis5WJvGKyH+dd0a1eMAOsPcbFSA/5BDrSW
QUcFcFQKU3AZYjbyDe9kn1E2wpTDFuaxzIFYmp4YrE3qw5LBRlIoeK2oCCmfkhQaGUVPNp/i23Mv
u67zlKUIvMXHvYQo6JqKgITnTbddBUqk4XMx1nCMQDxqrl4Gg8u34tAs6dWJjycLspE8mqa5h7Bf
jZMonBT1x5EmD0ubA/mt2YPBSpIKICXykjntErftFBWNWSzSIR5MBs9b5xOfnGe4d7QsuO2oeURk
duP07Pm8cagnFKS0G8huCc9Wxm1bQguBMSJGO3aIkkyNaO4hxfDdA7R8DDgAJUN21rzJJNrMd6oP
XaqOz5cor1atMd+5vsjFSauslvAAzQ0HJ+r9pkwNJqWw806T4zhnsWq4xc8qwpZG8/P27mDG2A0p
X8wzAMCSpGiM3DiFbS2R/rc9aQ6+ns03sotcCxDc0BGSyATcTOr/OMuBN14by4gODlKcPsAueJVM
7rwyXdr9I84N2v2ibFBeCpELc8kdSYMnUVEseWQO3RDz1dRl+aZJn3NYs76tN0T4Y2TQxPVVI2EK
GTDQqwqFInuX1odJAHObzK/DMfaDVsY3XxmRPQ0u0i9EHor9cjjxHJT9Dw4uwjuXbUASB/o+YeZf
46XRvTmLkO/Qne/B/Jx56ykYU4FSoNyGqjAY20wvcFPTHEFSMlsGvvLh1kyFlntQx3Ra+MoOolbG
1RvuMH7zJWUh04lN5GT0I8dCkIAjOJOf4EZBV8+4DJvrAPDYNr/1RyNviwsIv6pSoimfIQiMseIL
nOkXTdaAX+q5E4bvgwzr8G3Nvv0+mriT00kbG7E/CQHjzYreu5aYVobphejnW7O5nxSgccAE3lI3
ltH9pqTTAtwZcHJzVpghj+prNmsKKREcvH891x8RAKPxpWR81wgtwL+mxT976o5aNRK3oxSpnqCP
rfZR6YwCkCmvutHWdlwmzNxQasRHFIH7sVqY8MbRALaslEiSGGPCDu7blL88pFA1HYeKLGZ/GFRi
Lylv4zXb+KxFpEUFAGxpESEDdaOL7Eg5uvYBQi4I1R/ThvaEedbeJLE3nQMr2IpilyL1Ve6unclJ
pD0Ij7aAlFWWsT1FedSUvcgHJUpPgd9ylUTB9Kdy9kgTkqDm4deYSVZnTkEwSKupzx2bllaIg+Ft
c330IHxsp9mjJUHjqOPM1kHNE87eft5j9x/XB3FcEKpmcOZ9Uo0uC0xHsiQQ6bPNpo0dHP8+MYXo
7klx0Il3zrytBvwtdDRbttJnxbelicRgRSTqhB45blLMovmKBqFV95XRtNp0bJOf3Mup/euqd/UP
gXfsjWOt8v6D0b+hlwobuSxYy8dH3NdO03GJVMOHvcIvWYI5YFKdrSA4Q34OYPK+x2jVEKh6a4k9
Qh5CeFVOkI1hHHLs86Z77VrNKTBxkcqY/mTYj948lHRvLmwBJQZwdrQFqtAPCzJS/eHGY9YT2Occ
lBJMo56OTsGKN1dsw8D5o5dcPhwMGIeajix3s3Nt9z8qVZBx9YueuSoza5us0ueCechcbQZz8wcA
0cgqXhW7Epdjpqhpmk0SduNlXODAmWHsSQjLMVPUtQ4xaJFWqAh+hMnq/fblh7F+gV5Cl3X9Ws3d
+QoUPBhMauJBwfdkJv8+k5utITk22j2teB1GE47blXdkamaCXo4/t16pTfG2prTVMt/HRozkXyPa
v5ysL7YbbM9UAVbFngSqDEjjlYXVVEvWs43hOHY+u4vqYoiyTQtM9BlSRo+W7AB1f02LQDBGvTy3
ULdfsUQdQ/BZWsjLlI2TPzV9JLFqoEiN2Bu2KXNnhq+UnOWBDqzD0jv9FhH//uGf6DY6zYuSgjg9
0hSsSGifUfrlrOA62TubSXhNjzLFLruoJfj2MV8TNCfjvdx82QkC+nFd8G1sR5cgIpw3LeMsFxLi
9md+vG80LLVVSy0lK6e5AZa4P3+Ff69NJxeC8ubkq2xpCd7vS5YkfO0x9Jo0++08lxuYY4m4Jsm4
Pdfk9UTykAy7B1J/xYVCmyFR/+COgBHLFzI+bIHQ0x5SQ44m6oRi6+KRSNHZv0+1B291MoqevmGg
E+DXm3/ai8mj8GzTzXm/sT+BRxI10ZdwaFzYK/PF2dUJ9Q6pX5KJIzavnR5DJsABgA/lL8I9tr6B
4UoaJOR4d7nbtlqeAihX9r71ZU81heukkEI8uD/iO5AqWKyrOau4wB+fdGguB551Ul/M7dwURcZ/
dIyYva59k6jWc3g5zkZPi+GCBXdgMb2OJ/T6OxYPv42kXVsFL1RkvB61ki+RJnLoXZacTveWubEh
wNupfsza7oeKw3U2ZJDuYo/OMvrW4nvWRx/yB+pEQz2B011q8p67i2eC9R9z5T87bUFDWFJ+OJ2+
2f4DVwZ6pAchrD1EzDet8ui16u+aWReRB3R2soVsRHl1fOJnBOpaJUgxNmQvyxNHbsckqQxP5hrS
yHKVBAKbP4qKYP2RHCjhe9cwHXn8nUm9bsCoIKMrkRONjeMxBhPxlxx//QFz8B5BsnT3IfC7Ditx
Ei07A43/P75LXkH3C32J5DbdcqjrXctmRAcV8ZkhKsHAwgDVSHCs9yjsfwXKUmApdxz2MB+0bA+7
w4TQgwO5lnZh/T1hMYlucf/Z/LvfXbUk8akRYXtY2daP41k4BOBROTyzCKCG5bCEpumnF5LSafAa
wpidZkBClod3u9xsnvYsg2w4mlr/IS5vrX16KGWCoXbN1By5XatVOZo7oWtbnkEwsNp302fm4/Oj
MstMOuiSoJtXvHAOL3AvoU6g7ABd9U3SYpVz8ct7iKumUpNMG/FTgeZ3GbZzn6tCw0i/o2jX0ks4
i3wQGKuKZlHstIpovYoVbICX4T7X76/WQGh1i0mYpscepe+0RhVwfzudKltTFPQnCy7nzUtefzG6
5v1iGrZY4QtcBENWDjk0HL6FxTxhbuWr4+L2LyvG0FNYwXTUTpMVWErjydiK7RGXABf6v6XbYWqK
MoucpNN1dUwyHl82QC0PMuFPOlWc5qJ+c+TllZ5XBAQOIiFHXAXwUi5uZ4DqsEYu+VFf8jsJeHj9
hMefwmpx5O7KJ2x1wn/xGL9XmdjYUXnvBtcw52F/37T0GCY10sUPvuFtAVkrii75Qw/Mt03M9H75
WFpDsL339+ENMW3dSOVMArI0Z76mrCnbu0wzZ8eKjzmSr80IzHNbNz2QovyJ4usxjJO3QnE44PE0
X3A0gTQEzwr3kw8kCv88FfCgjizU1Nc22wwF67b9aGepkStxyUdATbBcE5jFmIVlNqsD9hfknS8n
adTbjn33IFvI58MODbC7UjZL9mbUAJt5ybxjMgnp8KEv7irOkq5y876Xr0vg/vSjX5jC/c7WXZ6O
cHKTCyckslVCtt+DYNP/oI/lDF0i731DwPqOduaRzLAseytWHXHChcYDz2AKa2UgVsg5j0gq5PKe
GLZJcz17TmrSF04s3ZBRjcvIiyB+Rz6KnoR09eMOQRz4oaXLlSP280WswgowjGzfWh+BeoF3XqGd
Le85pcabeXWt2MaVmOAOaE8i3UUxS2GyW8Kzh8DXh9MyAcAsC+tu+rdWcj8HkeZxqU577lKyLYBq
DBocyZCvr/eDu9iWKSGNi/A+WXcYROmgJnZVMHJxOi0jqaAf4k2NEhIge+wNXJ5AJcWROYkUMKNV
WmpEik8yCufD7i3GAlOziagLheN4qUuPTm03VbQSVRxEFv8JmRAbZLw48rLIpzXchVdU37rYq1r2
wyMtzeIpfD4FHcQR/aWouHG2WkORRSVDJ/iQCSuw364yjfzcOqIX/x+iow1Ft/eejPFWz540DO8z
OX5lNZbMXEBwhb93wiFK/uaJ7GWwZzZeqO+QCHiyVnbO7P+c24rKKHSxme/S6DpF4s7I8iUEhkIK
juAPHbAnym4RZsOeO40UsJUsFGsVCQXlVWDQBQTVHYLjP1LEeUfxbFlrvcPYMWicjBmlO8/rUGGd
6+/pL98mvgs8D8usqvrBmsOHM1jg3vQQYsQVrEEjD/vpK1vJNluHP8fu1wsAzy9K/r3g4KzGUhWt
OYgnBIAkSiJyqvkdXqHo7/cFn7c3ZK4lm5vSoP7MboYWxeycY4gorYzsEZKB0ioyJ+muvsmnf72w
Az7MaM5P/ll3KmSPE1bhyD8NB5TalOz+ihAWGXRTI4kamU/OfWjGUUlqyS6wP+XtBVAVybQQxcgB
cuZJW9haVV/SJ97YHJiEF6gLJCqqQQE8sGjtHNh4aQe+Ue2hXKADOaLCakZNfCwrjVHPGZT0rs1C
M9/yEaJ4+CNhoMuN1snZiz7t/0NtAuc/wipm4FMOZ9/vy+dY2T6gcv7BaEp+yT8Y5CpF+xdH/mN0
QGN6enG0JhM6JOV2YsETq+CPnTp/b1iA0fQFyC8bDp2SpDsO6Hmv6+7ZOBk8LHpcu+dfTEaHene0
/8v3Ipga1jiVuUT6isEd+P1nWPJrag8KHFOuQ0e2KP3KnYGuLTfVOA85eWVujn3hXaHbuTS/sQB/
42zbzlz3UJOua1T13jjm9Any8JFud4LsMvsM4FxRhHjE75pXdek1h/Or1vkVJnEZ7esxlkyKSVpX
K4Fa+wIFlXCVWib/k4eiKQChzbLKOSyKrplsNQGmTQNPObE9WmKS0j2QQNfQkkCW26Ar9F1Vgshv
+81zkjZft2+kNZQr1IjMuj5YyxcCLInrIcAL6I+TtoBSQM5gOYVzWWS6iGDrzpWwBXWYNvbIr7/F
2sr5TSi9+Q92cWH0LH/nHYW8rFa16Jwn68mXbLARg+ZbESDv4T2myF5B2oUBaHFR9RWD11sC8Kxd
7wuaelG45oXqAYBK2lipXtb8N6ybhSt3fBxwM7iaamyC2+LCyv5xJuAUr0z7wS+iXgYfNukXL+L7
+qlXOESaJpM+rsvrPY3uNSnJzML7Ci/dG6dWc1EOERrCUrFxTgd3whdabFUWHhrGCaCsPX+VUcCS
KK/d8+snVGXsAdwqWY/rt2+diGbvff+ewaCe+G8SY14bVZQgFEqwPROkyqPBR8Nm93OyK+/Rc56S
2kDVh1fc1MJdBtwP+HeIbFM7/ZfkCS3MCzKNuQElXk6kpHgMRaFqWbw0Ozm8d4QMimjEuc9kzF+n
7UfkdnmhI4AIPKkAogyOotJt5E+xtJOrO2ElyWrUgnhHF2w0C6ABhF0Nvr2TCBbiYbR1yDR1LaRq
3KU1MlNfqRgNaY7Kl/zhECXSaqVjNcdC2OQyLNxlo+QZxY3Bl+DF74N0krM/n7SJXero/CxmO57E
xBn03qsYj6gBZDXVOwxANXi2e0Rni3osfA9crje+UHMMDh4I8xP4QIPo1yQQZIVrGg0anLbVOQSi
PDbqmI2mQfhnJwJsBxgbUbWC2UhercJRBY52PJkT7aaUTCFqCuBouXQ66+pQavePUiu3ePBHZ5TF
jZzszcK7NnkUgrM0QBsPVmLEfacMycxCi+ofEsWmevS4WBo1Hrr0cf8hsH0qGw91eJu061vQnUA4
30d0ESOscUWjgsbvUnJCEtl6Bk3TxcPKlmFyZWzExV7RGfcrQrsFKmK8IjuHbVb7I6a/TFrujVpn
u/01GuTe32p0WpoEPSPBUukKN131ejL7yGJyEz8UZ80HFDg/4/su/LOraFY3TmSiTqcX7cLz/5cs
nggCUD1RAzB0PUjUacjyXCclCAmjjR+mSPFudSkkHN0eDnEBRjUFfPOjs9he0rGFeknd9HmypvL4
c9XaI7eTtyQVnF8d+uapigSNZihko6vg1BcKm+AaNVOeRJim0OPhCY/adfaDeM56LOnK0QEybclr
cmHwFGIKKNMa/PJxMnoDcVtMykAxd621ukcoBwsGPr5uGo0cQpWSXdGmVq5SdT5fo5YZhFaOzSzj
+wKMqqiccd02qJWynJT8ExR0sH+GoEViFSMdl+UzIp2drnGUiAO14q+JkxMvBaGW9okZB0BySEAQ
m2cHJS0/c1aAQr88+0bYEt6GDsWqZScBrYz2ZESjkgv4o91WDzS0zAaJkqAOZghSdCFdpFGGb6LP
aZZUn1+9dfPjpb/RFA53MU72/pusC3FYm+dQVnrEPX1Hmw4M72XtthbkIstmZW8H+vTbAyNe1yBH
ClHujHcnX/RRPAPkR7YAkJtYkcyJh19/l3AhZiyy9Y8Oc+YwTGOvJRMBEjO4lFj3a7XFadPxRcvl
Vi/LKL9J6mjjXiNJ8Idmk2glIeXM1cPf6q821K5L4zF1ERdQHSznDTl+G3GU1umeTo/jRvSDVKjn
Yhau5wkPzG1mcbkoYpesaNVrL7qibc4B/jw7eJK4vOHA3wfRSWgoNVzmVmfbDaNv5HlvS4mYI34y
Kr9JPQFslyBXGK7QMkjir2HKRjYsi2atHsiy6iiIcNc+NuJSTVq2qb7KFDjhMjQtwd8Y/8JmHc2/
4GOjjPRZPhzrhvojdhMtw98HFdh2n+QXNg8QmjB+BMRQKq++0emAuL71hzpQmKRf1e4yx+PZPaE6
Mwxv1zZHwOJ+R0nIpWOKGerszckC70LWD8VC1/ZJ8QRVOjnTz7wki7VbfYL9jvVE3owFJgqeZsoP
YH/P6j30F7I5Y5ICelQwR/50EY1dCuOw8fBwgDVmoZamyCx343qKsf6+0nOQSdfZgRLm1exy828I
8yJjtTl3SXKUbva9ejGUX436JlxJLmrF/NhbeNEePSSEXFiQS2Lsdfee5uECNC0HYcAnvoplLL+G
yFFXq0sCY54JdvTO14aLSLcdZCRtv1blAb3kQ/RKYPhbIy+bgch/yKN+0cjZeYewLDwGDJzBEDhX
coCr4a1i1HeW0gJajPKcS+6D8TpK5bk5Fnm3STseNkIv3ZsiBQFhFTJDNw+bHARxhr5hSK0kvIAG
jjP2mxvOKodRzWCDQYm6R4WiSKqH5CRcb0cjhOZW3ktpCj7TMuz7pkrgupSCxusQtz6zNWGPjFZo
yC2+96IZXpSpA/gKW5wCtJv7f9ZY81uakpvuJWIbs8UrcPCMOATR7wTufPip3RxDrym13I9vwTkP
wqOfIPM55xXRwfWtXTLTdMJG4oXrDO4hS4RpMn2IUaukgF7hW76Te0W4OMPSs17T9hH/ZNGXO/lc
UhE1mhqKQXklvE+BpMTAkYJVqd5UHmNIMZgIvgV3JRxReovz4YArE9IkpeekYiynkkc3z9Og8+Kb
MlOkp8oCjwACGBnUa8SLVSvimVP4hnDiNJ6QbigJPbdq7dcJNGotI8YgDYFZ66aanFrf1ToIMqxV
6RNAhIE3OnzNFibQyC0Pz7Bq2UkMA9NjWq4k3tyIdGAvnnFN2waiq6u8lHQ5ecNElCekFl9zqi4m
XDTTlOYLIqaFfMtchZaPTXkRLz1C0/xjy7r4seJ4l3kw9btozM+kYfQ6r7NF74NOARUT7wxlXykP
AaGApA2N76cwX4WBja2SqPb6+7WRIqo4gz6RV+lFNyK0kW7ipeF6s0vxZww6YNaEGIYO4uTkG2E4
VqliYibySMKK+SkD3joIpd9HMGbWGAXWr0++HAL/2YD/kolwu+RX32V6Soc4xJvaFsbhFjCMJfv5
DAY1+/M+jc57ycsL+1IfWIqmpvPR8OpxaEFPRibTpBO3mFfRpl06CPIQRnzedHhDPQScw8xmDT86
ZVET/mhn7DVWtUD9XpE7dv2FT1sw8v7SREmCAb4RE3MadMhBPbR2KCpjxP4RI6LBWcLfLDAv1ohZ
jKfsqxiVDal42q7cfenKVsHqim14YGbhKWjfo4jOkr71DXCzavXW9L90Z3fxVcmPjc+RbzvY56iR
UVa9bwnq76DpDez+ysqWCa+OjMKoHE86wQa0Ca9ydcTlxRsXCTV4U/4SiM4RLKAy7K+bIxZm0+sg
xgEfbf3l+WAktooj3u8DZJSi9TXWm/i5M0J07v6W6RPXnIp1WMVu07L005bfyIv4S3zyvxp0Jqrj
IjzlrPfPqQyRJ+I9fYgbi9kUErHGPnnRCSVewk8R5h0CweFlS7axl4jVkXXkWecS93bSDit0A2Mj
khVFm0ho9cPlCsIc/kSPESWEnibt5Rfs/CrwCvq28jixQzy6ecDPuS7inxKr9HpzlTB9Y0cSA6eJ
52h1D7yHf+NjRVjUpsFBAEDcZoPTFPk20fIApJor/noTi5odNd9MG/ObTb2XOwZ/FWwpN/tiNVx0
3eDd3S0U8OEH0MQ+PKcoaL1TOTdBe+3+E9ETG6SnF0nxRZCDypniTVwnEeqkyu0GOT2YGBElVpXS
9QGp6i2SXNNN7YQ82kgvuuyWBf/Bo8Foni2X21qDiMRGmGI5KvC1XtyOD4l3LfxgGAXYXzfO/Oll
7B4NCxVkAJAhW4ouzevvrR6+uvPs0QZQ3JXpgpC4GZK9qHRTpPz4QNLAXQyRRKrr5GNEi3dqJsCX
9io6m8kKxtPdWBQxlSutnZQS+V4tnOBZ9Trac6qMTUTu9wZvkKPkVJiq5gkgFZVIzFUI46LyfO8p
oT7KfXHUQtpM6pel/T/HmNb9ye+v5yYJU4Jtb0tFqZe8cTQXjztvaMGTAPW5Z1pA5YK0nfE+TTEL
52PUgg3FRnHeVvwT3qNpi684TPWCKUeMlYRPvOZPDTR77SgmH32EqkHu4bwz0E0UBzYkYvnCQfPG
GAU9dhggcnyDQE87UXjpwFlpOrlPGaMnn3JyaSETz+gzGgo7GjLMQyQQCN83Fv106/KSdkUbGKUH
LKdThjrl1uzCQUgH1xT93Go/2Cj6PHVOROUCxvkjTwM6iO6wj4iBxbC2ZyZTUlAgI6XpO5FeVE7T
IW/EHdIOMATomsHzY9+bOYlGWKWkpHV9sZgx3NcPSdllnZlNvuwRw+2aw43GPD8XEJBs6D2LLrR1
jOfw5E2c97Mr6SFbJ/8BmSbp2EUsivr2yezWzcCoFlDRtueYimH3dyuzz0KXtQIm0cTXjfGOwAKj
CUoeIiiWPo8/qn/ungkqxXd9eMT0ndxc9j1zoX4tTDdfu9QuQoz5jQuIvqc8CkNPTKrkmlvdqZWR
Hhr1QkHzavbq6WKMN4DRMk9DK4y7xNN8lO5eR9iRCd7VYPQA7HeIUVwEPQLhJf+TPNSnZyPov5rP
VSjfnWaeMTkebMD157hsA5sLy/r0DiNC11aK8pvS4qC1r+vJMUsqzSLag4r5ZyWd3mGTUvBHr6bq
qoyXRTLpRHUYqqEb3med0bwLLFYS69UPcwvJT+Zu3DgZj56hlBMV/1aW3jCFedtsB1uxkTv+YWvk
BslMEbu0YP+3kz5+qeutsvZuTtjKx9mg6SwDaFGdxyH0KQulSqFm/wpTAKkIf9C4UmY4DFBTh7KU
5zyfZm4dUPWjyXuQx0nadZIZbKjwNz35eoSHHll4WBWEJkyLmslBq6PAFusODdTFbwpV/SLNvRCH
r+BClhgG/3Zl5Edbmz+MvNC+7npy4gpDMnPh1OIrZciYOVT6oei5h7/tG0D+VCw5MQW+sT7vi+ee
YMP7xUGkL6OxgmqjRfa7e0T6hm3UfHabt1leoR7kj82qr9Y+AAd6SYqgr7Mr8aO9Wvjib/Py/9La
oorYfjA+2mLqvD27eO9mvYzR5uGrbzu7sy7dU1RvsIqGCFcWlUQWEhKc+gqnF+2CiH8mY6gMPWxW
GpTMwQZUJ+n/BQVfHV4dHPtPnDhPmzycX+lUXw4QTf9LQyj+bMVnHMWuc/rpS/J/y+qKRo7oj2t5
7LbG5RdwX9gsBRCgGRS+DiQEk2f/yodA3yM55MrEetJaioKKJo2Dj4TeYeVxDC0+CR6idtGMaa/r
suRRnJ7lJ3odJGiw4K33WPVsBM0+tntQ0g5mNBhGqZgID5hmgVvL9GnGiL0hNFLuLZ85zV2+AahV
A3anE6ldyEKxjp13EA0Gc8xbj0Vv+oBXH6qvcbh+mFCasLw9V9CAQwd1swXiuGrTVZH4s7Z5QOgZ
I0yjDL7z49a5bMYvObE2PkuP+B/5N73g+GIGw1by/b+XvPNk9KHsiWhW6tOl/iTvsQygrYVzgAQU
PPHmtgpAj9UzpKzJEQwuygUMFUWM9GsIXpOrFUAoRtkiEpyb8CnLvn2kcBKItVXYGY6KWKsYQMf4
gqRu5ca9vTeoiW7cblEZJkNuO7pw4ATj0XC3Ix7NnTVXM7dR//rXvTmLHhuB0f023edcyOwwq5jp
zrQTted/I2iif08BwocS9BgRq29vP08Rge3JaZLCh7cNfp/jFec+NAmE7yzzD2J8Hn3umpFdlsuB
XD99E+x1VEJI5jAJAMPeke7kC2caaAc74qinuVDbw/dXbsrlqug95Nndgp90DjQC1qQjNaNSnYsy
ORE1Nf9vIzwtuf8bg0APU0msxHTLHOwWgeg47MwDEEWrebDjoSbCjmye6XtFLndP2ErBt6dtgEYd
NXN50Q7fa6fi6xpPN2qiLtNvE++fMe84JqZP6tr9Rx8N50iiVCJEikYG9Y3aAIVCsLto3Ii15UP6
5kIgef0cQBzR4+td9umtKORcQ0BV/vXvqDWXP4QwYafcmNiEwXhHEC55Khrhq/xoubRF1pewmW02
Wu6TIcQCzDdd7NAn1xYEJ44a+f7Oium/pXJ2oWbOw0EWHwiCJJzDVgBXwG5LlJRikbAgUO/U0sVS
ipkCCjnOSiOiMzu0nxjT/9pMsgIMGDRVG0xd3s7XatdzsLYwXZQb4elvV4qZGvMWUIWkmzUo6CqD
WICg9KvpAGrn6u6B03M6y7UCnIxTU3b1GwYdjsH4HPzrRDULcI7GCkgwxGhDlCsY7+zxjqMMP4jB
LKT4gE8rBJBB1AzVh2MyZCGKDrrs/JcOr3V7rP6Z4KNgDBV91H87HkRZiiioIM7hh/LIjRFgxgR+
I8QWdmzKoEO5T2bG3iuG9Wtv5f1PhqUbV/UfwJ8kKnvSn0aVNW0ScFKsodbDazhw/AVYsWe8WUdD
fNDuUGn6yhJ6um+Rid5I5pBphwk2vQBSniSr6VqsylgVUMzeaZsmK6CWXikjwjUwZSwud/cuAE/j
XgGLZImKZ3/EwsuB94OnHrAGbVzzkI2a3Cz3Yx5bBE+BmM4KpHe0k23hoN3Ntd1Z+4rYvfCs6vWo
4retq/1u2SI36sQNwuM/m4IeWzcWo0brC+MH87N4iI/T3NpK/NDrhQ6x66W8q1kul5aSnMu/COAy
Ku1gdie8vsSlP1KWH1F/LKwRZ3T/AYRSqZ1mAz+p+emeAeVQv7xYqKemvDHZjMG85wjsWTUaH+So
qkM0ZDvU2zYoQl1FHqE3pUmvoBbEzKvsK0rUULYiwVWBdb9fgxmCJ9B3umCa1ZIoGEebx/yrMxdv
sjk0Vt/63YJ2MsXvlGdazruzSXpuIAmF+TAPoaQ8SPdgtVDFOEwYhv3ahhd6AAvsDO5IVKsoAe6I
gml+ktEFWcYH0SFb881J5AKf87wEmqFQxDkIVIt+QZO/M7b8ODsbMUOqAVv12OxKvC+xfsKvLqpk
jl3oCPE8hmDTKdHM1LhSYsU6EiH1RaQOmKpLrLaKGDc9rPpN7msG86678hN4hx4qYNpoTZQ6BB5S
Kwh9JMUZ7TeBv4otlF7XmWAeN7LEROOQ8d9ebyhs/lNzW9tgIPKqn8YpNij80YsfwO2m9MarJu4c
qWuUnXVKM7JlNtiOsybMAOTb1MtsUHbQ5bfcMyxQL/+auHkwHbItU3Eex/YyjsVDA1bs2VLlGg+a
EWEgf5i+i23LeKOrFAOKEF6ctBsobW9//5udaz8wE43bN8C94fnmtm4pWFXAfVQwkvWCmmVtsMrx
BNh8jMDCnnzkTOzDgP4h2Tdi02ET9DJ9QcYppMk2OVWJvQ0xQm3t3Olhhn8w2PxMCzer1GyBv8pa
+qFyTLjBqePH/39LVM1VnZsYbv3vr1/ULsd2lNC3AS6WTWW3x/KLDysbALOAsueg3gSUpCKHn++g
rPEDbI31qKSPdcgN3vK8j6D9csg6RdCL1Dmh3lZqjI63HLM3lr2BUSgaldmI58Egp4v/VOXa6el3
T0gXQ23UYKJ2Wahu6gjNtccF2uxqFfY5GfXzTsxlPIyX0eQCqjPOM+4sivo5dOlVRBmfhzyAnwyX
EN9a2X8+VZn0rGy3+bxVT9bnzhRH7qVzWa4DADr2uNmkeIEAt6eW6VkxmAVrxoj3zjrObGlbFbXh
rbH+n5H270FyrnjMdUt7xJOInovllH9FseSjB45NJkZIp1/J9YC+5vN3/JT6sY0nnJ+yIqtx2R2W
+N8fsegefRymIAexBGNpfU+ykpwlFOVFc2mrzs1juLBeY5tsQBCOfCu59dHwVtV3QzmMF6OiKpIL
KV/mZz6g9a0g9AwVxlOYXLgMugl3XNmq+ToxWSb2rbLnttva0YfdLlxygFh4Kisdx9gxD/6s5I1i
rwut3ApFOS8nSU+iO9EHXQ7MptVfmXrbC6hFFlJ4TqEvVVVEG9hnd76t7dH40gNpfCscitrfU2P6
Z7RyASjxMDsgab8euzp26HiLvOgwW+OiLyKyYvD7oQSM9Ngk6e2dYunlCmEu8iRwnpcFR7pXc7v1
n6PpoZumkiodjmqBTWA2AVWIPcXaCzIYZcBVPBXWINIJOZpY0pD7jpy0nDs4IFwTMcZ8TN9l4pXb
jNXzp0GiNognA2WYOwi4/VOq0cPJ5KupnLtyYVBPERfhtzrHR+r8G4Ys310pywOD5IPH/k8W4chW
OJTQGBom7w7SWfz5MCRnQHZ8DRBxstlnonuchDqrPh8s8IiyuTFAdxzjdmrGI3pzll8TDNaoN07b
ft2GXN/LKWlChDOpF9U3ICFBYPjjK15NiA84dZdxPTCvXMzw1tIU3F22vW6IIWKuvqzfZRI6C4OD
25wxpI3uW8Ef0DwYL8mgki1W6ocMDuuzRgJuHc4JD1pI66CN1FCt+tNw6EbDzuIVsoXrgGSnddCc
FEpAu1jIzpyH1pzWBfCWY27ex8z8ZUfCfw0t2ikt2Bp8xNgjxGRL+Nco58ozNn/TyvnlKZ5mDNnW
9fnwwZWx/JjWKpWg9GPxtMQYQS/ez0beMANzmjhIBzmiQev41DUrfGKmZ5i9ryhHYhbSPE9m96ck
Dld1bXG198F/UUVWLby9EC/xaWMAbPqSxchx/ygDMk9lFYY8QRLZf8/NEePKu2x9i4dvYhJ1Vn+x
UGzb+03PnYT4DGsWrgLM2uovbQ6FNl670TtxYnbb4UyMbHdVHnDOv4qmy3zjriNkb1pHzK0+tOZy
Q4ECz9GMhkemX6Pg4BMuugbTJBjQPBoykFxBnJE/Gu5anmk2AIieUM/Qysk11P9S1WATbmGUSX0Y
ENY4T/rLaHue4BzGSf6tqYevEQiihunmZpGSmanuVT7kJ8z326fXydyok6/zRvVZyD0CVLYAF6qA
wMTsVmXTwU9N9yKx49lF6MtyDRtkEg11XRYIK8fLrsc+WaXsmwq/ZsBh7ibcQbolfDjmZwZfN9Ao
JS66CIzIUDV2jDGeHObEqGK2FubRSiPtMTBUp4YS30xE6wrQxRXKwGutAUurvKo3qKunVGCXzbbi
UKvwmJP3q5zNEru0PMb1ckRs2IERKw2Bc9z1Yp3/eYtQQ8m2H7DQRU9sMaIXpmkxPBHFrE7Yd/MT
PNASzI4XkM0Gb1J4FcIT2oHzdCkWmypaZpsVx/iegCCN5Ve0u93uNU7he4L7tYi3tZuroyf5czPp
fV9dGnqQ4YI/1ofH5Z4puBUlSYilvCl3XzyVDakrPI/AkGxjklJdNh5tM1ILr+TBoHQsb/8gXreU
424Lo4tYj7w/5ueGSY/6/3e7Nuv3Bnm2g6qzknVFyZKZrm7rvASR3vGs+26LhxnNBhfKk8fr54KE
DCJuFOjI6zIMrM+G2LpaZIvetMBkMwsXaqclEyna0MUDFhPSLpUPISdsrU23M948sDIk97l8cGO6
Wd8uwL6kD5GnrSsRuZFUQk1lNQ5HKJVhs3SA/emqJ77RSin/jJgZlmZomnP+STKelXCYYXbVljeB
+H0jOgaeBBYzFsoiHpXUvIEX1lfugUQ/DIHttNm41pNQ3JXJz1gUl4IFeLD+YQNpQdSZOTesHyxE
Dzyordfw3djyBKxLsH6z+KumAxTtkm6RR7TFDyiLXi3xVIGZGzwo3kUA8nzkx0VGq9NvPlZncPVJ
fsny8EAThyspv2/9YjV4aZOansf6xDcwRF8rcjhCPmPoiHrRBpoyxeIta+5MCEzZc7rkG7F1Ae8y
8Mrn0G8CqDeOfB6g4n0ps8EFrWW+ZYT8BEfsFBtdNRiZPuhepMEn/8Jp0ARHnIhuXojwpw3jK8el
5M267S+HN1itPrEPQrzia3q+k5vE5rHAYfMleU8l79dNsZTYFIC91qb/lbivqIqcEi/y9kwIyl9c
iKQCMqIWbBSFfVwfJ6nRlZwcCzYYiFFYRbCEmMyG560TNUjUZzK+jk//9fSWPcKJ7Es+XqA32n3U
w87vBYu9G6vvwL3TLD+dBKeA+HveE82rbLZOf1JVt3XLoGQlzoea7Vw01Klo716GC2Z/U3D9LYGJ
IIXJ48Q2XvaNIb38DUYkRsYrDDjpTMpZn88mdR1QoF9i5MB1MNavG6XLzEyNY9znptUVW13WDY78
RvgZvBVRCCnDf6/wPKrdFGenMvcNSbCRmGwzD9OE+KBnBlv7f+ROfkZHuxZQwew+REyOi6VBDyVh
uEb/azlzqBjGUJh2H36xFdhkoc9Mk3DYgXJV/r+6qJInsYQ3hSDhsgxcU2R6ByyJ6trm3k1hwCMR
2bk/FZhJXzrjqSwMa7WpFWD3jo2vuDPcoqW0S7eoG5Rt5QVPkg5pGGGfbrLK9FZbjvqcvYDnYa6/
n/fXE0NqAkagGhAxVI2iV/QRZwXnVbcAg+3tNQlZ4aD49ofj9PBOApihcjHwYzqm1lHUvLF77TIe
MY+8+nIBxy0JQ3Ap4os/VMzKDXZBYzHRAtYjvzrXhBYfWkJpr62ljDeW8cA3pO0cnlWulxOBmSVP
B8chALBa2KcNn61OGEWZDekSHe5Ud85mmDivC1DAFAi8+SurgH2Nr3/Xyqr5wNXWW0snrhBXKtf4
fjwBmLZnS/jJZtMDSOfX9b6AvVuVXiG7MT6H0CB2dPqNwy7ZESencgAJOc0tQuFJQx1uQ3w6+4tS
K935hGtEnCAlzBdP1t0zEzPU4lSNu+4bPxFefDWLgG4NYBMumlOmlMQgYN11jHAdpfxnNFchVw6n
NY8rAbtQWLzOHGIHzWgsTVwBbqTx73OIQnnVmp3+TB1nlMChpnxfGVMMqlrtd2XA+jHMnuM27fAJ
I+gLTsdHVR4XID/75OT9lQfG9YoArpyKWTreM7fY+KeinrsOReNVatraF9YHsIt4GoqBhz4zKR40
xqVar5zr/OTgWTt2wImnNS/C29VKAIDi2DZMc4ryKAOJYQMRzS+Up6i1fwRI7CAo0xwQoYXvQ9Gg
qeBebXYL6BLG538/c2zqeUcojH9EmV01P51b6P3MGkXLB8rvvKSy2C5GKgKv326K/Sek4kB4kh/y
zlnM75cTp9gO1UVBxZq5Gbf4AQmTCwWW84HB+go4LiyC/oUxb81vMCH9hgJrT7vTw/q/XsiUoDR4
OZJTIzWKfVqFmiRT2O/3DNAH+JyWNcAWir9ojNGCG3Yb55klAQvauIb+IG4UsYFZGhM/EfVbAKHs
UNsV2PjtR2za3uz0+F1RYrqhKG+FGMoyAsgy7pYwn+cR3fg+ysc9pceD9wUD/yLIxPlau5b34KXq
y9dOkEX1X9/Ey2FnT7nRQydAKx4coYQe4Fi39W9tIcaPlQAjQJ37orTYQD6lVybS7zEsOEVRvo4C
v7L9dVgYkbSRsv61CUjCP20/N7Xj8q+m8rM6p+gKNew0keMTeSKI6SIc870oGgv1EhD80xWUC2V4
+j5Y7Fb1UdrzRdoeTzztzb4qAyXARkptY0xYL4b32R9qCLEW5YyOUA0+ZuTgzpuGvFk8XWSKXDIs
/d9DIkM0yi/4PaTIbbK3h5V2w5prPQl73JBgt0ujBXu7DMoQ4xxdhXbUymK7GNcdhtmo07amvzzb
mNiN2PvlTylYKzmadUP4F2t5QsK3aV6vb42+lEo8KQa+M/uhVy6dxTOgu2dlny6SLitAJiEeFn/e
ydcdONC6dqY+5mdwS3WrYHuK2XdD2RTvqYh4Xfk6CRQ6RT2nBmk7QoCeQ27meffn2pUcNXT+Flfh
afgu6A2OXDuUHzGuTqTj6OGu+8U1t8xxP48dIwBNfkPSEUwjHP4+1l3s58rbpRvtlyrYFAnDa6T/
6pGQWvTtc5uvZNTQjVEYUcisasH1hbajpnzvF8gjMtlwR++JFx7ktv0GHl8wwqXueWNpJCZ7eoJZ
KRee+DoJ2SZ5ACqvwL6xZVaSfkGkeAjD6ZbOsOYMeC1gvCrGAQAF+akzct793HlBd/e4rLuXyWVM
JiH0o88h+uxt1gTFmP1gIG6znoq5ArRRy28yoIz2Oo+6hPykWY0WcVTp4VYijwBbDqWR/jNCE6dz
zR7Aw+GYdbrEZxzuE+GNTkkX1qRs1M/8UABsxK1Ltocm/fe4HsLJyC0DBQ9iOxu6HIV01A9JYr1r
zn4+gCLxVN/pZc0XQ2WN30aSprbastbK9Qzk5nwT+32GW3RJ8VdSeZcaEmXKWAtk9Xt5MVZuFVbI
Y1YrJ8FIAevdacJ7dOprQBeyNrDzbnf4+vqe3V4U0XVuiaIA/Q3QwGUDKsjA2sVppfsdMUCOImuZ
c5kDuyrbnwFIE0O8gTlVcLklFSaiqx/ApfjaBWUoMQBQdywsonWrYl4arHLbbNi9ZRoqlZ/X2bUQ
b/X4CSaHBJPldchIn1nx4QvXsPPdKw+U6NtUf2s5gtlR7DYGRD5tYkZHt6/hc4AeI8MxBQz1B42p
AaTUuiuGTBztC/D16SLXE/qZklSdvHbC2MapWuxWcgq6WU08T2djjHtUXoh5qrmYemc7Oz6xK4Pi
e6EAhkTeAhuDQoP1m4eNFtzIStB/SS+EWWzhdj1ML0drtHgKhLi6hBX9ynPrhYAIP3VGSc1yCSuz
wkgFPqmZal0j6sspceZZf4KsBMEtQ95SwvPmnT5u2Z/pwFMIGYWF9l6gHX07CsCgiRF6NUPkyRG8
pvo70v5Y+V5sLi0oqzJDH3VbS4VNCSTfx/4Lvv7XCyVQo+mEiN7CAXrX5IgdvLI/Ml7yE5YtYz0e
+/GJz3hb11RFgb/VrsiXCoX+ZCZCb2V0rUmlLzSWJzQgFJjIsTRmABnNAUoZ+mT0GDiidfPQyyJp
5cl6weRyLGILJsaXzbOISRsUZ0qK+t8Ibblz1ZMLYTNZDU+DGj9NHLfJk2McuqeJc0OKLDixviF5
w5dtMcV/mhcR7ShOUxcCMOdGvT6WX7MLSzIl0PRSVa3H09u9/w0gJ+cbwW6EP+dZvS8CJV2CXbl9
DSsQEifW6LbTOltecoZHLEL5y5MZiZrcQOGNrpbpFJ8xN2MrRJl1CJpiT87msDKOA9+4u5Sterbb
NqqySUnaBTc5AYydPBcI7Lq4AqQhJRmME8E0rJbjesIOzx5d8z3U932nwqYmCWA6ee2TNDFpaLwN
YY3f7zzjBn5FfX6hu1m8DJdZTp4VV7bufb16mVQtzb91RfRZTn1+6fyT3GQfzxHbApMeG23GvRpM
zGneAO2fcsJHsUPtfDsRzs0Y+ep6XveOA958nX4b2qG0JnlVIYCpHCAw62VSxwQlICDns+szeDr7
1lsxJhp6Ceo4k9nq1AMakASfpHatD50Yaw3bfIUl8tFq2U6ti8gfGPKZyEbNFjM4qdi3EMj4R2eK
obOFJ0xeksbd8vAC2FfKx6g5oeoko7H8p3zsJCeJLVS64DhXkSjgAz8Zt1mFZviRP7U0f1qhh0GR
9dqlt6ffQ9ZtUCNxmnmAdOwjN7smEKIrywPZWGpcVcmgyZJaKIOGhi9hTclU2XEMsp8kdgimVTdK
YH1Qp5SCWJWw55gVVReqLGcT3TIhHA7ZlElK42xc+otZslcV0mv/hkq4l/ZlU6ReiVJ3ESJapkSt
jYfuHvKLfsFcMyJ20TSuvobgAKKbMWWwEdy38M8gXBlbwGI3UuemRr5mXv1ylwuN93YNX0NJLEJG
lUzOxEL/LafIocJyOXyBYKbJmeq/7aAp8WCfjtQh5SD7lZeJQJDmmF8WPvMC2YTNJTXGd5wrsnjW
qNwesacrAXYvhGMxbWaYYYJzIIaalh7q4w+03XLPKAKUweGxh2zlF6cXgsx42MUBHtGF41jIRVC6
/R8RbCxQhPJGBSDbTnUR6VZmAwuXE/YFbtvvxmhHXCxY5RsYLRzbRZ3l11KJ7NGh5b0foihySbq2
c+w7pYAagQf7cwfpKN+wr/Gwmzp5vrf9U0SZEx1yG24addoIjBmfnWOfDmGlsAnIyu1Pt/mGxBdz
O1ZPsjnZnDUuIY2UC9Di8eLTs71R0gYQPLSSS7V918/BbAB7r61AJeRo+UcKwX4FzQ8Dds2N7Igl
B1flmf0yx+FNr7wjZXa74bBI5D6QVc7PZ001eYyKwf/xZoZUCVWi9ZyipqE09H4gW1rFIM6Rl0Y5
dIB4e38E2F4RQwGsLGRjsvymPMzvCvuldtsEFOytt0eoPnxIKopc5Jg51E9G+S6KJwDous08tWI0
h9xuU9e8dMcbhu9aBIaGywPy79dcs74EnsiPpKlmU/1TkpEthbr/s37uRst5lhj3ptNo4gyxrcVS
IRHk3cDMzE6hsTJoxIqUdJ7TIsF5P9IXnWUF97LTG36eRwT+87f8b+A5nb17TI2Hr++GJz8K/Vbj
+/3h2Db6Qsm0JfpkW84hvEsZ4OVEqigitVX+ErmyW+84TJ1psIrwjRJYFn/HORQusmXyFPbsXI5n
Jr1CjzOeL7ETYRdDJ2N0Z/XXxGFagHbqKUJHzgTEnwJlOZ64dF6IN8KUDA/qSkfpXjqLVhCh97+J
waFdwVP1AmR4WrZxh+Pl5nrfUNQBQzSojf361sK2aXbYcXA4PdaoLCnQTRj87Q7MoNqjSFjSpI5Y
dMo2bhEdrBFFho35rqDrQvTm/tvgmQ0lbJ546bUpy0uUjoJQyFy71mDKg8saupyB5LbuSOZ/sXdJ
9o4qD76h1fkNcHTYTQuCReAKWf080w3qFUluakMHeqD9+8IP1gmjuZPCqAV6SA/yx/S+m7caM54o
JFym+UNRcCH1YitD8CawjZuJ5mqLBL5lbEZjrgc8MsCb8/kfnG61LOjzUmIk/UVlqk85uTg6UgVW
8aW6RBc3coBVe0v6/Vh37j16zEeKR7zDr7G0Jj6YG4ADxZUZ8cAGn83I0pfHyMYw7eY1oA4AXtg/
u8XvT4dis/jH1MCu37LzAs3uWO+LcxDmWuV2AkTiWShAVxE+pZbNVb2U7C1PXV/HPCkRLuYAvRWJ
e4ujSKG0vsNlUoEVIZrRPKwDuECQqp2ZgwjTqQAlY6ooFCP7YwQh3bC/aaRyuTsaS/wsc9Xx2RgY
TA2cKZMLo2BpSJIPgsTLxQbqBGCXv9WjBruP3skmHeryfCBiIxKeubuWjZwWETbvwR5cSAUG+5zC
CGZ0w/aJ/AkJG0i1mrRtDNMJoSE2G7AzTr1RK+fYjOEXnER4zwnJaHAzY0Bb4Bgglb2bOIV58HUK
igYU354rUiAKlHYP/Pg/A/OW83Vr72vcghagEZZnUZGEhMsYaYj4TfJAKplyUWguso0l4HRXy0E2
bFdMOn7UkuUM4FBqEagYyvZnOb8T1+ObMvlISII5gRWgMONni3wOQke3l6l0ruSsZJCI+9hfROwH
D302+MlRbazYTs+e7SjyvOnO+fjkCzQH+YA8JEyBi1ryNbcjVBhjWETZU8Y4rQUC3g/+nP8q0+wS
fCAQMK3iBBw/+H1qTswxcNEDHsTyMlKTD9sLOXBG7EoSVrhuFIIgzouX3O+nbuMsD1BLK7ZAmDwn
8fzIC1pk+6zL7kLCJiuh3s0Jc66HQ4qTDgDfzGD1gTkBJc/vuXb+ZH0rfTqAnM+Wm8HdSNmp58vN
fvTo9bcCbsqDjnBmiSDLcDWGBZkCF7R0rquGBxcVgo145dbsTv5INBnk8TVWxjI86dDqMJG0fc01
Gu2oOe4a828ETJRSFQqHvvagQSLyqjpSkoWLDZRYfCfO6SzPau/ps176V8isX/h81y5hBSxmlqbO
yIOD3rwHzOs6kD2MJrYtmSkbj0Lq4R7r9GIMEkOhzwgC6TAPLSelSCKqEYyofY+HvHPtPe33KeHM
5Wd5sTNLn04OmNBDDz9PKz5nwOjyubdGmy18z3QOQC4YcUszEtlZ7yGtdmU9BsilVB1v9NE4OfM2
dhNVEjUq2Qegmsdgd7P83FqpwoenEol+65okITcjp6GtzsbK9LroOBFqE77oJJrBmCWeePs+mV8j
/8IeD4bym0ugr8iD6cEHGgfrYgXOXrXGfns41K1rn0DxBL31hAp4JfdhUCEbtugPgtPEZExMTjkE
jyluuY0sSwfNFOu2J39e9SW/r18RxYcddqMiKA3yI2oJrXgXCLNIpOigtTwiK2UG9d8HAKZ1pICf
dw5d3ksARpFQR65sBNIcH1XGX6wbfZGwU7CNFUIan8Krd5pyqrQQg43I44rY83ypVsJrA/bseL7m
Fwyn1hfxVHkxNi7CozvZv6HKx2xJG140dWT0qcIbP7nz2azQTAQjKQ4CD56zG7QwoFaYmD+kmoOo
E2tBC+s/cmTGtUoVF3ZuUZN6yL7ui2Fzzpz1AeV37dmCbINpZcxxz4lXETv4uToTK5ay/QGtsN2P
QHS6qpVZIp8ilp3xZCVUJrKV/bMSUyuqQzTRlQWQyRoY9gLA2v4oHdrIvbdEC9aKgrAvuJi/gbdI
peNRwOWKUAqjIbN84B2gz/LfHylh9Oy81wqQkSxaYSBIirZNcB73kkc6GFUWPUY84I+gRT7nReTu
p8EpMuu/Gkm+sDXUwxQEAF2e6Ael6qXXFcUI2TAo60zjRWQ8SsWgovkXuZp2cTVeaF+VTrB/bVM0
zv+aWmqG1su/pYIfjaT56bDuvcqPOY+B5Pj7iMLG0gzH8NatraLBwLxKkCTiGzqZyeY33vmXhkgY
0VrPPL/u3sBdlnlanfqR7JZsU/3mhcIjYdZcxxuP2Foons91JxepQUzDSmJKtIkD36eQlYLwFKgU
lI68XDf/WROs/HUdZu3O2Yd8248B1k14OTzEjFeQ3QmHNlRzkRdaXycMT3m7JjLxNqY5yt1oNy2l
8efNXokkLlCtKsq0gwTolXOSnqWFelq0d/RuQo6RIEvXS6PL3jOQLJNAxALhpj5UtbnCWGVCgqzI
zndFStwsgt4yx7Odm0j0z8HRCAASh2OcPR2+6rtPA17nuaGgfPNgpO1CSRc1XziupvmDctzsiHcU
ugjS/qiSbiP24lS8KeoiSebLljvnY4xvCvcYbsU2ZZofh4/h1Eyahl9RlPVCQJ/dLS7nYFzb/31o
+bdBN6QVeorqYdLJBN3Oe1Fpt4tZOigm8Mye9UkoGgPsqdU3YiUa0ndJQGvNHfIldpSkLKWnGhKF
T/GhLVftsXlFuk5OvQMkWtRU80lWaACgL+UDvlx2PXgoXMmfFnZH9R8BH9CEZ7DOHdgfJn+HOBx5
dFgt63JzrMy0IlWZoUlMaSZEPgIdeZCMiQrllSeNQi54E9AzBQEAWNxPjXkNtLch1IVCQ9KaPtjZ
M3P3qY57VnoKhpR5Ts4ZxqE16CTtK6yP/jI5crS6hm7MMIXQhMOBp+NQIEKBNtxlOlgiyI/xfYI3
dECLaH8PJpMwA72GpxA1w5TUuz9LxmomaFA6ctMyL3EtcpmE4qMiNL/odFG2g9OPIRKF8tUbBdKF
0CNnCXYKHlwpFtFmkX76q7IylSp93WuoAN4+yVfKUIKoL29GislrBXDc30rWFpkTXn4SKKKEoToJ
pBDllSSXCGF/doIXB8xQ37erzIsOhR/i4EeOgNmg28pQCT8/DzzsN8cvdH5/qK97EIoOGiY64200
an4aicKtdc0ObKscC6KOb1rIPT6A+mmbTA+gdNxCGRFZyyRW/dxGMtka7T4UMOUxc4G/BiLGpvPx
3fWOj+mInH0IlBQr1IZIAWdsdbTaIVYIonrx00vJquqRBhbPSv1jlD28kAPUVzHlwALoQdrxish9
13tvt9AbF42UutSmNYDl386c1mgYwaxQYpkTbE/9IaBx2UFQTQcQL1A9TEkDbyfqlMARqdjKKLaf
TEvxkx03IYtsuoCTmSwg9kUXRoqp0lbEghGqNxIGVLgtgv0EqtxTmb/j+BNCMsGEu8RcrNmgZvgz
MagRP0VB1XfVqgiXVoCkEcrBEarv0+c2yHBlCzeU+OSE5PpoJo/IsJjmq7H2oWy2XjiV+WGuDqYm
CZ2Q3r1F3NaL3LxID+pQHYZOzKHA0eJ5y5Akkce5JFlj4RtjFJM//CapXqS4qGJOy3gg12sFDN01
qg0/Hlyec+TC1Z8iE7HSTKNPax8mHOfoneSwLi1gVW12HJanrfjS0B1kdIgHzsUalaLj/1MH5yrx
vb4C5FzRR+BoWGwna6Dt1x/FzsbkjZj0fI2CnxJGtYKcCozRc5/IUEC8v/cKD7MAoqf/m1tQM9q2
GOdE97pqo5xl8JjCeqaj9OnYyolE9TzrGENZzCQ08aMop1yClz3dvQwFI+LN+JQYlMzKKaSdVpuR
ELCuzxon1Ip6D1ShDJa+qU/zu28HMWGjUEOSz5BIPzoOlIjpCfr5g0X0DHtLrk1gMFfRHBvTM7C7
DILVCX4QcEi+/OVukvhhc4EVlxd4XZRU+nbrk7A0CsJfrdxHBK7xJlicvTcJ2RIJ1Wujh0neyGU9
NniHd/ZL4Pd/lWIOGy0SuM9wt0mARguRNEKuRhvt27dqfcIu7aW9iRqmjQGZQlPcwkaErPB2CUvJ
Vod/uhqggHzJC3v2p44OQiPpOiLRiW8ZZlp6cnFwPdph7g108oZ20fzs+6IYCrll3JAO50YJrm/Q
9Chz4EyCnCFFygxghtaEB4x2k0r0kE+7OjHp5IwwGdkgEWHrnCxI71BMy5lZBLYNK85wIn8OlrQG
VJ263Er/MheZtf13+Lv7onbW5BhW5EGpHAIKCYJUFYzAygkOcbjACZOLbNQQlLMmSQn4P80FKAH1
Kcuj+LNxbiGUqIkxQ7EvAHftgH14zjOCUXqRih3rvVrDX24JAm++sGzq81LOqLksL+vICeS5gB7U
XewCRa1f93y9RXDVPVZdiwyVJc+7DlhFi16r2SYIIjgNtCPcczYL03o1eVvEpQ07eDiSOmgcZJ1N
lMQ51HWrVoklyswQqUJFDoRmRcamejR3vuyjghKUDYS5y6DL2jyloDDeycVAur8umYrC2afPWt+h
5I9QijUT1k/wz8mJ+SzTVN2ENLw8Cge9VftXxTf6ZktKObNtFBlygXEGtc54ZR7kwRE4CNBf9mVv
3xlhwkdVMJfPNGtx/3vCXEx6zNTi+xvmh9ol2uMKBnZ60SXL592094r5QEbxgFPAy5TVFAkJsUqL
y/DdpPho4AD8dL8IaV3hZ1m6D9w9xrCZhBBwfis2H6yq+yDY6X7U9PhU7wsrV3poOjR7ZQSWv4st
bmEE9+I3S/A2C5LgE250I5pUgfUa64wQJY+ikpkTysMezPktsNPVLZ9gKemk5+57qLYDqTkEZFkR
8ETgHC6AzNbIVNIeRrYIZEgH5Howy0JP0+MJFJgpK30MPUvdxHfLo9F1xsRdHwAKOG08Y2ZnUDu6
GMIcL3oCWi40tR7SPEI/WJ4MRTsVapQx3c/zPDccdbL8E0oUtMlvRoTP5p/UArmGc2ri2sHgnPf1
ktnFjLvV6f9ggep4/hh1B6hULpSc+36k14MUzhhBx7FAeAbgJaHSdrmZtTE4OZXk76RVjnevSBhC
yXuznkvXIV+4BiGKKBPWqfF3Sj8h/XYDsKd5qwCVtO5w/+H0HliMam5VGtgXBciGASEn+RMvaZuh
Ow8ftgU1IzjDgdOos+mCXIBm2RhVa8/N70xOQgeyBZtl59lJorPWTaTXbXt4bqVc2E6BU45paG6A
/+NRQJaS5SVRXMrR5e4EQlNI4H9Caw/8xRso59svByhWiUUV/vSh0g/sVVjvIshF09XwwwGRXhg+
K485y7G8NjekqMCWVdxOzDjBKbAcHGDxHD9s6TZe40u+4+vTiKl7usT9pfeotXpHErholoyzKXGh
F4Uk3i7yiNpx46hDWxLxViSSfpUjZCYDm7bxPVacLTn8hI1x+uT+azQHrzsQxTFhA4xYk41mNA79
2xoFjLNXEv1ggdSb46fSufP86qeGwZ9BrYfES67eiP2wvdyqn4ch61rT0Pqg0rur/igMDbbgmf87
lNAyDcjJ2sk5Es2rDDAjHtSKtaOP+bBDv0QwdGImF2Lw7YxNPPC0iiua3JYRMUD3+CCZgmJTNYAs
4Y5ZAwCBZsKWAg2E3OJfF+H6gD5L6uyvclKQzvtfLhNwakoV5BUix2fkV33EyT80+WbQJR8qlQ9S
ysrS+Wd7JCK3W7nAFzTtFvEyUvbC44mGJkrHLxRboDYOCEq2wOwBhmd7XxkmEpUdMZ83MARNgRAw
Htd+WWvy3tsLzk4ng1csQCS3OBOF9lVKXvW34ZqOGgq2HRpDxchcbfV5VVdoA0YXbhtUJ9wa8AYW
C6akTGSzCNTWUuw83iNsgk9RWxGhRVONUwES7Kyzmgzf9YpD8IxXTmtrqXbaOZ8Sz7X3Het8/dZ1
0cFr/hwVmmozn1e5uNYfLOpgIIlBmuKi5VhlzJR444KKnVUVJXu/vhOWOCNKttDGaH8eTNi+I8Qr
etc05upCt/F1vne7+dN4XdIAR/98GcvFQSqk2RnOWGgjoGytWVy3DqZvKVtPt5tJhKzvNvhMDzHk
ufypX6yk8C7n0h4QK6DuHvfRGaDNIK6C7D3MGqrpKQLWPMbWwRfyyk9++ferfpKpsdVkjjO1LY1X
iCVc5jE9nXeiEy0NSWwdqkhZjj0e5rA4KcttJ+ph/E2XRlASiLys4x9l5VXnySY7oCELBQ3osC1T
Y+e2mFbCQCWtxuLrupkZL1mH+/4v3EsHK2adDadaFKHjaxkO+8fTqG1TYQhhEg5pKmR0OakTOOSD
mQe61nxEE9c1skr80URn/D/m+IVt/iav7hZCFYEP6fbCsygIcFzI/VhDzps0OnxBHUXr3sSZSdl7
G6lYjrW/sr00+axwpfTaAUSRFvsiqmx4nWbDKaWDcJK2hR/9ZRSC6rYVHmjQKfuRZGdStHsS4zFk
t2+bGgFRyWb82ut+7y/2/ZofJCE7O8KipT/9cknI9VIJHsnIlC2jjLDwmBuTkhq8WOZC5nHvsLVB
VbXwMnGTFg2x6Yh1+dJbQogYvc4KqdsI+inCrh8VwL4S31SMTuVZIIFJ7x4eucAwe5ZGWplujREI
U3oUo1yeHRIOLkEbaxLsKnXJrlDHsngooVEaN1SBs/Y8o/woR4rnKOtJzsLruZDSAtMec3EZGd+D
Jra7NDvN2tuujGqyr0JRsJdvmLipFUodOcg/cdMR9m+oxW2fourGE+YSRdDdCNJAm1Bds3bqZsF7
fJXT+H1ZxfA0w7f4Ug34LHD2UX5RGMBSkVvOX0tMsunYz4LEe/VoF8fzAN27cymOiw+D5pZOHbt1
jEPpTJseYhPEOJj+ea0KGLHkr7s76sCG3HtRLgg3+fvsorZNPL5dwMko8HaiATcpzOKYuw1p9f1m
l2rUOQIhSWuUR/CbBVptfWGSVmXaLLDLcwuJqAtjYzT6gH8C62FvhgkGB5EKuSowMO+UEK6vpu1k
I8M+yY1ixPDnN7bkAbD8otlSE05r8sfOK+dZ2PMgmwpkH9H3rtkrXfsnLwNIw8yaaZqNIPp5Iqua
+nXNeFiCnOBWlJKGW/vvdqQyIJ3DbMyLcI53ncsSz9F6D0pMN5k2/QuICShXkjNluptIMA2rmBsA
xnUHXvXgOPlHDvImdrUgGvFj+JQ5mMVTMh2O8aH6XiqjuOtgqEXfGN6heyIXqfKSg2wi47YMHEju
2wm33bFAEBThxx7mYFj/8eF4I1HRI7t35i/BSbGCosQIortevus6GWMpn/Goda11e02MMH17Gb6J
G6PzqII/UFK087esGkEyV3AcsUWg5NHikXIhxL6eNPVjxGeeZr29MuRYJQmvOPxTFYLanhYN+L83
liTMZK0g3A32botnvdYkIMiSL9UUnWqqCWbYSm7sXMlVmuwcjABODjCE66dE4aFpoKPw5jUEaFdE
eP9/SUzohOKiY3ZWIAM/yL7ZZbmInSVlDWoSmIsdHbqWOoWz9jWYb5bwfboUZ0YxFXualgHejWGM
cAYI0tZeFGbTO2dtBiqYGsOfSJBEjL3JHHVi4Pvf371/AW9b2JYPzLTbb3VwibfTvtVOc8ob3rcN
8nIcZQFPE88IYwQ9O0MaRejTNA5kF8XsxytvFlkH/h0/GXYSJ35AFmq+GAkap31RNWxDMpQuB1vN
i/BqvlVRmPc9cDv+KT0pB2ZNvhG+gXWvWTEW1Zr+OeMk1f5bAZH6YUdiQhxaTEt66NUiLnNUHLfF
CwCCmtnTDNVuBSmbFiISNa2pq207GTZKTtXk9hfjPF92YesGZjvuStpCGZrEKyEV0D5Y2IZ7VKVp
7Fu6qmIGy0c5fa8OYAcr/XBQWXiihL+yoovdMxNZg2U/3qGLeR29lKh9YFPrJbRsUFFWlsmGvu8N
4bLXbQRcoxkOJTOWvNw8/1NMtr76l+zf21Qh5g2aFjwNmJmAtTKhR+a0THkrzRanwl18YHjHKnZ0
sp/y9gaaVoDXBWcAPz76+jRJQSzz95B4LwN2RpGF2MM3z+YN5FJfwtJrbA7dawB3ZABC4oAXC94T
/TiPRnzzVvu8fkrFCLGcKYYXO9DUYvveZs/YYcz1qRdgSpBFH2JF0TYsnQEA8yPUj4S40JCiQxrP
G8ud237lq4jhIhcspAMsepVX+37kZxL/0iijcCtoQF8WVvKR0GbuFE6ZjnVAlJx2NZjq4DCOj7LC
GLom6ztjeOsCaT9C8F0TeiZ9nSTLCAr94TGZ7JGwIPLI5GtgXF7Yl5Eqho2FLTd78WV21MLAeazq
uANguhoCSDZfCZet1WuPwk9d4p/oUvbkT19co3Em9Yn8hZdod2AECZpVejZyLrn0GpXm1iFZ9LE6
LCsVwqKogI5n3avRMGJYGet5TdbCrrYE8WYVaYV6JFHVP+wSly8WENmwwp7owa4lnfwRDkG8zkpZ
y9n03X97OQwZdtlQxyQxsGTcFa3k3/0uI/3Rqi3qkE5zxtIZR+SIG+JgECSTPtgKtSacN1OuoyPE
preQCfEtIsSPGMSlhnkkRoodyFYjqbv7HNyQD0JXfaK/050s/J3HiJCPlBWa7b0Mg6TOEZ7tKsZ6
sqX9OIP2IQ7TpmnvJoyfkC27zOjXLdI+eHkpgjFI+3qOhVZn6qG8jHLaBcpJwThvqvhAtRcladtF
Oq+qtSypiRRRsH5sWSpdXXdOATR1Xz4MzUpwiSoKDaqgI1EAxH6hCLcsRRVjKFQe3MMuZM/X9Iiy
BudEuWCE2e45M6WnyH6WW+9JkCHZgi6ev3vWLvnC5fo8E7pNouyapdw5zSKaDUvXGWLqd0V3OIvF
ZHj7uXALbSztqMrPreKVtwqxlqY/7T7RXFUx13V2JvF/3SYS4wu4BJXr5kcPKU8WydKjCBNtqoC0
k1s5+8fkd6LDprh/8NwBRSQI7QgECLcSrsJsAsmQb6ZhxuYGoPzWpICdv0YLFKRUVtX2DaoRQKv5
5xD3YPi8HL0R0q5RLIfWTMJwyD+qYP2d4efUu0M0N65znCRI5WkSi113sR+Id9xGbWAawaRzDs1b
Mvcgu1NCbGuNuucqowsjVvsJP8HqerB0R73KCcVpYm01p8Upqtz0It6UkKI6sgwDf/De++auOMKr
lPdsg7VgZruA5j5QEXfdwHNd/Wx8TDADzhg/OUh9dnBUTcJB6Ah/0ox4t3d7WedNOJH2aXoZ9MOJ
1qP3NoV8nwihU+wZDH6NZXv5Rcpp2ilVzxxi6q/SYEff855wMQgif/Amwz2t3OR2ZxE6YbUmrUJ5
z90jgbkzfyiyDsrKn2YEKyWasTkSEpCgfjs/Hso+s3UVYIsv4dud2lTWbb5NIpU3SwI9pwxMDLzS
RGwAuMmyE26Cs0IE7yAhoZQblVjd9ZTpDV53mJc9Q5szNdx5+xXqWUnLgWEUGelU/YB4wjCu9xkx
76zgt7sfpVYbPQqJnJxlxoxnh9rkxrjpiRw5fETer+8eFBl2K3C0t8iKmtPMzcUs0SGdq6JwYYia
odeCsTbZJHR1DuzGEC8xAyPKP99uOuLu1CSoiS3B6w79j2/5l6rLfOeXOgO+EQsZH+/nVFRAeQ3P
/GVKozFmzdhXtKUxRMOOjdMDaRH4g4nwCccDhUYjp1lin4LXE4DdrqjD7YBtQG1Kj8BZUnUbmFjr
G21qe/hDdP2Vn4f6oI8u7zFn7nw7QVzr00PK3mghNwakNDZMEIWXP6ineG/okxkc6kYJaheToOS5
OA4hxR5q5hSCmwKCUNHJCuVADeGSg1xGkqiFyFpH8CmQNbSLdGMmQHiqkI7LQs+u+f151lY931R9
H40QdE3qUoQjtjU6VqJo6gOz/1Hr1RuFqQiN+KzTNPA5W7pDXa9v+X/zGqBG0a1MF426ldOlBxdc
PAGvcIucKdlOiGGeUrLIY0iVBjvo5GgWfMOlGntc2E+qVZ0ZZZWFfYuR9LtqNCGQPH3tK4/6ldZC
baemH38i78Ody0F/wRO+33Gh05RFirj2xkqy9T0w/TAvyVqwkYC9nj77NTJDPiQmIwcYBOLQAChz
8L7XxnhkWMNC7AGFk7+tNpd9EIN9AdghKnQ1DVx0n3Sfva1u5QjHFdkmJALMwE4o+HzjKcepxsrd
UJFk8pJYgcLldEQRWI0a2c1VOodib0MO07s7Sy6X94Ce7oELbyd3id2f0IG2OQweJGX2TQax8I2F
uzrpwKTPtpj5iu7QzfZQccRu7tNd/VeGShAvNa+CdBIMsC2IBK7UOk/0T+nWYiN9kvPuUPqurtd2
A/fT/37OlyXKT8gt1p5YtarZvGz8nG6sZ4JErhg96rMpZAW8OQsZWztphDVQwvoqF/xfCTEPJaUv
4wx6lI2cWRn2iOzMDk0akbq6ipc20OjxJ3JFvKNwRnHUhjKGjz5A3keryjG+LYyEb2aKo1VrORuA
e6YpkAvB6KOsOSqJThnB3HgjwZRr5mcHPjdm4exKrzBNgfTyKA/xtNwhkX1a6wjrx+KR8HMar2XV
fNiNrlHZ71/Bv4n357jYUhVZUcWG9tLXVS9iG9dshikEXIndpn2twIF5lQuVZOhKAEk4WGx8Y0xi
ObtQhzY/CfYvDj8tdf4RBtHpDRiu4DDyy+7B+jmGnvrm4JvvLZBJMoHGHTvfzh+909exzO2eXeGW
DZ1FlTHDxTm9M6vFDmpmQshlIJVkpZUt0WI3OHUVAqRkOGN4rz8QCEdyxNU1VdRh5rodF63rQOib
e+zgn87A8h8ackkyhbUKBzvDUVdY4qDpNUMBtkshGKF8jxcvWPxPXILSUg3BC8Y5PdLVgbFjjiUr
a695qpc+xlHBZSl5wTbAsb5LDRIxS/fv3KO57dKg1m+xrZy7zSI/QjugzZrQanIaH/agbPv2bkKr
CU7WFNTo3XcETXptXHbm4MyeRZahVVPfHqfaomFpKLEOaO6zdecROswlXxUMQGcqLruY2L3QfBx3
iTigO0EH51Fj2i+nv0kouQlyBIJPy4Wq+M/6VEFn4yJ9nbnO9y0v5rwKFBvYB8IY32qpYI4Rs6ne
d40H2DRMO5iwIJ/LH9pbSe4xoloP02thp5B1IDQoqblX+qdthxAXragnDMNm8R4N61k9RGPvOP0k
y+KBJ5WkdOJ1xrwu3X+RY14wJ/BFPMrqe+AQHWBOC5nw9AL8QY+PMDfCuTKy+AgfUgXBfnSuk9PK
pSm6OubEee9K/Pjzt3HNHUqSovuChCUrYxh2CDRMkFusJ4Vz0JvKTmPnJV8wOHkf44lVD2K+ExSe
OFfZ404By2vZEXif8bzAEha8yGSsI2+DV2lBclXyejogn+ujuP0flw5FfvQ6RvL9TPOrpAPEwB/x
pwkdMRnepkuLfAG5qmjul9EUhsYqrz0DqXlqarJRg9swaVpi2BqiBqyRIVMDQ1tBr7b5Jf0O9P07
idshp7VtrVPMjFpNxUEz7nSrhy2DM4vmU8YXAHndFFRnnYQvJYNVRP+yGxhOT+C4mrRhrgCHQeMt
qWvS23rM3pOWvXVx78ix94MZbImRMcGMk5D2Cq1L0RbHu6nDmsQhoJ0+ubEF6uUz2tjHedZB8Ky6
rXQjrSFmX/BWLknRvGqB/R9eYCDu/S7rOYKN1Bv3fkDCPHTQ1m1db4P87nGxmdIrxAnSjU1SDPm6
j6zuy1223FJ1S75Vk44MTWB1FyXRfe3YxnG2Ggw+E0jqikdO5sD7pFDL7vrnygz0hlFjqF7WPegB
aFIVxDAOCJJtsap+y11fBFzoNvEipWTskvGz5C2jyUCe2y7AXe4D+oOjY3qIpVUBWHg5JEdyjcqK
JBvzReVVW85vwHqudtv85xyeESHnR6r2xKyN/TDtdEWv/woqpN0Jd8AkPp1MYrBMXuQVE/sWdlrI
36vTqUJ0C5IFoxxA9adPfadt6S2RdDFTfzeZU52gLZXanW9cBw/FXZlTaFuqPX8wBAZjz6BDlo2L
kryp4UcRefaCOYDEADOzbXIyB2EOeed1YXPdgHE7CjwvmzpfWwYSUtWpaxeRCAETS59mE/dKHEqg
chPjZEDs+1ayhWXtGxZmBE6td86eLyB/N9mrB2LquncloiEjAneSHcWiyBg41FQu+QoraYXjQR7e
Go6EsDGoBmvTUTMl72RHzeXZdDFOGPgISDCVKFNmf7Bvvt2LV0WJDK9dBnpLMHOY7HLCAoQEpNQG
P/fW34uQq+Rj1n6wGnR5Ec6JVbSW5OAsapZm5q2zERRaV6+u5llaKagW88+3Fr9TEVrGZ8P2Uy+Y
8bOinXaXzIQH+Thm7BKC8VKhnbGRQws3eUvb/jGO1Oj3fWNT7hDdcCNK7Jm8GrIalfT+TW3Xgi50
Nvbi7cpZMqnTgMgstyspR5O/HWrCQ7AB9PD8U0xILXQxbCu4fq58DblFzyTcok24nSHc9mEFFpxO
70wZI/JvoVJLYfyJj1IQ7J5FCSCeHUk2rJIaYn56jK5FtEaX7K9bG52SahinN0y4DYyhgnqoM/o6
Ov0v4LlePQX2BpeYsK7xaSY6rNtOzjYBEaYmaksCdbMwYmvPTMZyFtUEy7DJ3+mvw7Y455af8Y5t
Get78V09kSflaOrTfxzgadrY90sGA/dRbwwmQPHs8d0lJWf6GnkNwu+RCWXRNDmZmZLtVTAQkAsZ
Hx4mPg8vooiVOrX0IFunquZk5UMrLsmFIxksF9oGXfjHXTVrcyuPWFssovKDtEuT3ZM4HPFNDVJK
T2xHxEdQ4PC/yIL3Cbattk56Z7x+RqXz007RPbeUQNWSRam9k0z7U966FAJmmc9EMwFH42Igx1L7
52ND+Gab1c0YbrKPXfX0EIGzNV6oAHAKTTxzkF25aIDx4HE+AXDExPsH/Y9I26PYnfASIfzRD5d2
txGqZ2cDcjTnREOPwuTLb2YptKwnF7hhIQaksMD7WuLn3hlpfwki3gjhjpSudGFL6SJFTSRAc5Yd
wXrqckcqpZYvUbKuUNTMjNyy3kjRm0hxuGrpA3npcLjIoSLqrcEolZfLpLDbgd7LNqmk+WhjiO1I
XgCBjyc7CYGdm3p5OhY77YxbOo1kUOkw6bVs7R8VFjM/rIjEJgejR0D8c8/0BP8AFLw+w+IETNv9
wSF6Ml5MA4hu7+JkwpPxL+ELSv8fc4uApHMWkj1ZtRvdCkRMKZT1D/WmH62oIS06eVhE0WOuFi7F
S2cIAaD6ti8n/Eil0rIRtIbhtab8+EzeAD3bNbgfyPf1zegYftuWvHv8XgmoIZVkTtDyjld7N9Pc
1iQ4UleLAHI3IK03InHECl3+AYK402pYKXIwmd/Qu5gsNlj8GVtQSGhUiI1VCYU50TYHxWXgnNQ5
glaHfP8+pX+aB92Izw+TeuDBx4w4goO923Z/y2EUz3IM0N8f8K2FluznoTzFXgJ63GFFOP1/2GcO
IYOZbZzSU01rXp6fs9MJg8Op1UUKwl5F2oVBzs0nDxt57ZLdp/KrmjxfpyqdBE2exKwIZ6FsRTFs
CCC7fd6jitOENIhgOUoRSvF367pHhLR7CTE0KkUrZKy8zvUEsGj62z9ACq8q9mdA6Cz5RL7vaRMM
t+rkSfXuAl6izrSRXxtSvQqXkKpBrjj3VpaVguYem9PdmYqdIC8frcfF16GRxfv5j+ZfjcKZuv1G
/QbqTr1WqC8efR2Zj7r9+h/Zgr+dyXXw/R1lXsMJXD6Ofm4mKHp28WeecGh4X2ZcH6fk+FZ0Xoj/
L4j5SPoKwAv6gpH5sjU2LlTpHRxeb+PwM2M7HBksa2nWyDOjfdGXUXOw4eFN7H7oEw7zQ/g0jdMe
fGxXmBKjGQMqAUTEpX4WQWdtUodeeA89MNSuEC2PLL2duPS80pCX6tOgtQqKGJ8iuphQhXC1FPCi
tq6raMHhTr3F8DJKIoIm0F/bPsl9fJ1GeuU1cE+9IVdddFL14GhUlK6neVl38HoBuBD3ZwUQ+MsQ
bMduxTRlVQq7eWGCvsijZkMu2Yrs7NQgM3H9W3veDliMSIOGxP0xh2XkxHGDBDBiLICVteaENy1U
BBhKZkyV3KHlGLEvVD6W5pT+XPvSnRLBvgrnGU+tVqDnDSnYU45BwWYlIkbkml96Jsrfy+RulYFA
AbDcUpc68PaL9nfNEpQMr2B2tu9UsAXlb0cMhp+nAUqi+8tpoMp2g0zP0K5YRIsQss8v9SofwTqx
+RX8L36v/wYBynIw8RjploG60PMnJqVqqWZFyuIVcijZ7Qtoy4HmSEEJsnXmAU75hY3U7u5UWde5
bx+7EFj1/kmUwHW+G2ea50bmcFwjtaYJEwydPOybZdPyeA5X7Kea+hk+MXCjxuZZz4LNhytYezcD
pQj7NiLB6QZxxzaLZskuFNP35KsRYZvZ0R4NL8wfsjHgn04FhyYwHAyepDFWxsYFvQb6XDfLW/x0
0N8cFPmvOuzMhO/5v5HDJ/iZTvxGJSEJOn6RD0hwZ0KZWYrOX43sPcdvI8rQHSXF/svQzkXnow8d
5Uj+uWl3STt4c0u4RmVnYusmFzDfSHQQMWauqWBp8KwFhCLTUczuKmH4s1RMNbmkp/2VUvHJEQ2z
TSb3k8QUqrDFqVecgwr1jf1YBfWJKmuB7n+Y7gjQ3yFERf5Rs8KsvWg1KeDyS0Y0MCxbWzs1IeZL
QpAdhd3e/SDmbXQld13TN1JLk8b/c7SgN/KEgPb6sIUpkhzdgC26ta0oeyaPiXxdx48pC4oE2MQb
XAICCaCjajBXbA7Cv0z1bUSyE/tMTqOv/vuJL+WIG85MWOSYznn9fGXmIJcEPBHeHToMKwR/YCu8
jyp+tNuk8pYze4M9BZlWV0hNbiEbY3kbNBKhCKxFEXRq3eZAG6nO4uruVK7gDzKdPS7xmnJRskH+
9RqJaxzFvNG4FHYiBy/aV9Rwfr+yw47nSX5n//AnJkEnA/7R89ykibqhhqWTZcJKJdYOOmx4vseb
QoR3n8ZNSJXnSJJTEb9iyBBCf1XAPOTeXeSveGxN+3WV51cGXglQB2MI9drSBru4P55mQ8ksfDSu
/NEHMWm1xULWxoKtR+rfTQpBQiOeecUWURG3IkuWlyBRvrSbxwnh8MFB4Foan7OCFXzHf+kNN1RI
fpgykn7qw51Pgx+rAi5ICGchtnaLuFO8rKnLiuHfI8x003qDjjZ4Huj6JKJE12vRdhYpGgrqDygt
pBTu+yCieIoI5FNSUgR5KwhzVeiqUhu0R0njJNA6FQHS1aDVuBxG/neKo4tsBpeiZ0LnPtKCqiGF
TObul3+vUgsiVyBTZJMhEtVlhSA+VzSJz6wpOPmPxmk3Zdi2bihJiFXwTdPO0UqOidwmlODtb0fb
ZlHWTreejcCKTBYhLqBg4X/Fhf+vuDj6hhDU5z3bwj2AgMf3Bqbuq4RWxQdfdbAfRqhJGiTfAymX
4y9W9McEtepB1LL5C3ssU05hdQC0kxGDdk2LLN3vmPHYFpfcbxJVW/LCNJXeB8lrlj7PJ9SRhN0Q
DD5waONV4O59fXl1s2DoUkowJlBU8y6ElHAEQBUXVVJBzr1o2RaQQZHF8wecdjCfGvhsVsX5z/yv
ATSYGSUBsCN/kRpJF2ORcxU1BShuJ0DsARIE5rlImXXYYTcYdgm8i8kCG9ncKtMQzWuvL6e6Iu8S
yb7LVzNtv8EEEDaQJpM9pZzp63pzDXOyQ8qtYXzmkF1mMWMuEZ6yxJ6vf8DHMoBm9PDBhRMzWAPY
UuCLZe7LO/tBRkXc0SW2PWg6AAM51rIRbVY5sN5syhLyM+j4x/veVV82t6DQ7B+bPnZ52dsaIipw
bPQy1fDqh0aXaRDiKdhZffrvX0iK8/1ysB/SmvLCVLG8cp4XAz6WSoX6TJOCw/s+CMY7prwuXz3N
NaUohgmbJ86/wIzzwM111oS4TZBAJaqy8WlUSWzVAzurqd76zYuhKgnWouS2AgAFyQ+UH1yp3KqJ
QVCHI8L31/om8NsMFpWvuCI6m1A73XU39ctq8GNpqRSw+jgt+Cx9LXzF0KcT8PKnY+RdL/UyE9/T
YYhNUPGqBle6IPethzNaWbSBxcmMCBWcUI/EstgIUMUBCcG2B7AJj6LzPF/UPtd99KaWwNj81Tyc
A/7h2VTW79zR8FoAfZmsUeXTRkb4pLMCs2tYM/fqJiDW+38j32B1Kt1GyoYy7hiSRrVZ9y/w18Up
6/UHMQv5/Fti0Nfo/VaSkCist99ajxn/8JP2sOVTA+xYc/LHbuPHeObqL1ixui9if5HB6B2SBu8d
KgWI9SMvoiL6eEiEb5a9rGw/cLMc4rl1jpJd2cuzsXhpEFe4cLPOWKOAdN8rDF2sk1e+ieslxQPv
GqMF685BlPPAXtNMKY4GgI24wHO4zNmSJW/uNvf5T57AWH1mDOh4ZLTEWMRbBmNSlgMeDYga4WqV
4hXiKDkKNKYbPSJelFvJc1Rv+UdK5FLlWR4xfrRIbXznSISXufQ6o5AQAYNR06izyDP1Kmczaqej
aImCNWy70mbJXLvO1uabJO6lK8K8kH3nixlrJTlaIW40broOZe2aivvyq015jFfbONQ4ffLHuOC3
tbupjXlNESfGxNgbH0GinotWVZCyxWyd2gpDv1Pe0pRaH9mH9dBkI5h39ansko9Kl9T0ZT6Vn3FT
e5JzjIugk0TcUPT7DLnubCuzhQ4CVangKaC/QmPzBhEuBa3UrWkkyGYFDmUPdFQ97zOpHXjc6zxX
0ZPap6/vgfOGzKjAOB5d9oeC1lY0IdhB6XKz7HJgBGOMxH6JWLmF+/cfvLEKAIOOL0Jmc6Vfp00C
J2t1XGpDEMuObQig6+HOYGVcSXkQpaZHSuJVOvsx4V+K7T7hPpTLW6wUMQp3B+4f34sLM5fJHpT7
dHn68RJjm+se8ZwYeb8yc2apO1Jp16OeIaH1rrH1tXFmFdpxfxuXtuFtVMBknZmPXiP9i3en5nVE
BpjjX8UjmQKgI4gtrkNoiEfhritgPPAYlfMk+xZPvcmw8uA5KsDjajKPb4cpSOhXylEmnFo2lyDY
Ny11rJ5b9ETF1TAxOQY+9X0TkrxuUCgtyWHh8WYsqmMJ1s192gUYsBN0r+U/EO+RCkeuYvxeVCym
Q+vjVrjRUWixD7XA8yeWQ5cyqdVXEHC9dIyY5NWWbai1v1DS+k8YEIv1s1vn0cpA4nArg863So1s
neWQA4J8cYCubxosZUBX+plwK7uxvaPE2Ygay2Hc7ZDAhaN9R1Rvsi4gC0GGopVukuW5Hqr8feE5
0/9JT/Ew12Yp+CV57Kp3YhqGmplb44BOFqJx4y2etSTgipHDlF+6MEzOnc/xWzMjCbDxnatSCU1k
unmsSn51F0SbSjRKJnPxLR5DhXiLSbhn5NizQ35qaxRnTuxZyzpNYLe3E3SXjsttYAqbPOI4cpUx
NZAJu0+aAPmDPTURwW0Cn9eQgs7r6gbXc/cxYEqqPa5tbfE68O3dACbU+eMsZE3suUkcul6nIDaP
JZKDP/83WtBd2rSjvVYZ1M4zJQ/vLfdu1FvnvsQz5GmDRJcBF6a1kvkwaPSFZtr9o4QLy05BVz87
rcb+D4+ZcCKXOyPnQoDHLS++ahWypllYeuoy+o/SFLh7ELg1VKou64b4WNe4KayAlZcM9Ve8hpk6
DJaQQAumxpURggt3hctp8oR/dpG+1G42sO/yj4rQd52/fZ/TW4SzRev0dg2+QYRCQKYmrGnfN4jq
d1zJJ9QQ2cy0vXtZnCaDj2utTDheCgGofQU+vFbbpWipDC6NUhHiMewBUXagzl29nqIeTLS3MP65
+aST/81f1qr7eaadK2ANH2JfSrViqg3CqOfcFCfrcXH0ZmSO1jZSdHWcjJUvjh+TLN/RC5Crsmvv
kCsymmF94F3W0qTPGX71W4Iadb7pdy9rxFRCWznx6Y6CqQ0JY4DKx5xcKFoIpOOr7MBuxDgWAp1N
qTn6iW3usNObmiu5XlPmsQy9rDjAXklP1Ng0XoT74D0LptzGrkxLiFDusTFWF1gqYHcHeM/zeshY
h/93ZAksQYUHdpi64LbfNKQqwZuKctJzzHDCZJB3qZcKi7C1eirMEn3WILMEc5DhE0dTpW/kplbu
zhLnplpj9w5fghWVYKi0mDQISCYhPLVQn2kLOxCqxbmsr1jMQ7amJJFIvARcYELX8EEbRU9OrODO
1GWA/zQNKVFGHsb0HjiIvgZObtgJyzUedwU6aRfW/5j1l5/rbyFy5aY1QLoC+75dA43rgccbAiHv
WiLmE9E5qqIXEW1t7Pm3fYALVLau6widnP2m9K94WycgSAwraZ+sG7IRDqD4a4b8IrstChxBxyCW
OQjo3HVOiyRKZVhKKxUPr18U/EgOvl8Nj/uMVpPGvaW9mB1rS0iszNg9ccdINgF9fOhPnnH8hPJ8
nwg8Iw5SblEkDA9+/WWId59FRuY4JCAkwTAbq1W34RmlGwnTtq8bMwvfDSp5Y2Oe6mltZk2tctXs
tnxCfpOONJZD3teaMVtk9khyJFDFXkEFOd0JbRSMxOxAPGTfGtA8BUpeKKud9HYCOmiBcC69qbdl
8xomo57vnBJdhbEbQzQLOZF2FkIh8np9L4JQ7KH4Gy6F8uoiVJhVYHO13U/0L2g/i3hDXOJ4ull+
+SUvdANhtDXblNmffaz0opMg9+xF2oL79Z1Q55rVh+0ldBPbdme+9KlcQ+ZBYCumnIXU9j/S9VJ4
8YFVRmME/OqiBgx3O/LK4D6q+zB5jTVPqH8ecJNdOG8kt+tXFHGU6YPN07yiBkMdOaD8H+74LvQK
58PLgZ5tIaDNlYvCg89iwf58jDkyiXRNaM6LW4Hk0ElRdODXy7njoy6mizgcKfqTY0MG+qvTBos/
Uj1PY/0+ZOVeCe3mUaq7EWYmNugydalZjSehT0jzWnidIxNyF5xcpz/+/DIOeX3nKrqztosTa0gH
tXbDpj9tojYn7YNk4bfKDfK3EE351p4P0RQiyppGwlp7rL69ACILtF8z7OqBQ2QE0p/YBFkABC8Z
xBsqWrnuYBA4s49BLvKoRAdDUANmmYK5YIFG21Wq812WzA8WUhPPWR8yXByak/4oP4X1cQTTbsA+
5tx9eVNxTxVYGN0jPwpI62b+JTWNA2SIXRq9kXTzR/nsSvCqZHchQZW+Q7Of6YmEYhVzzJDZBShI
RRCxfR3+TdZtxcu8IijqxtL7kcdxaWQsvWy64N21INLkMeJBv9yRhLaaJaZ33/Sn1ZneC9wGZ/dV
436Gr7H1dZMXFM+EnVcBAk/jCgGj/nMZkZaKuK5URurf46CaQAs9fvO8zDCBqT7bgOPTJ1FCbtMs
H+N0jOdH+c4dtLRjhF5y7LpYXKAzm2PngskxqJEkJS1M29287GyaJh4d/FYc/F6ws8pnWzsJ216s
cfpvBvi60j4sBKrXLaqNf0U5dooGteTREN+QOvDnWDhlWqywxZEZceERl5YaX29LfGQDZWw8N9UL
IuVxpiwy4jyIfqLQlVVNPvKbLbiX5I8g/3oVCQc/5MmGMDFRht5aWmZfO0FQ4OiejDzbxMcgJdSX
BJ7TwslRrU9Ws7x3OuLjwe1VzP7ihcALJ7XFcY/NtO4VgkZhyp3JJSSM4YqB8Ho2E0cqx0SwnybV
Wv66hfczPQ/DCa+cG4/dZwCWAuQXgOcnGizgxCosKHOEPygnjouGnVtkeVCuE5js3Ft1aY65BeDG
8kzV1ODqN0OXyHvUVK17E5KZfuvGxRT8joBcG43DXXVvN9NVAweDohtQGy3J+7gY2TNejCtlIeIe
N0LvhjQGDwu+66DF+6n1fI8aT9rfDBa4sjvx9tuCduGZ5CMmTKKqjMTJwpZ9I66y6tycdknmpryJ
yT9se4arD4JWaoREzL+ie3kQWImaenZc7iRSkroLZ+MQQ5dF0E2McGuQj8N2h+hQb6Wn1BhL4jzX
GUOAOUPE7jNsFvq8oEhJBLwhXq7pHLVRGJ00iIOIxF3op697gblSoCMhSk26PumLI7EFTZpze8jg
0zA5vm9ggYpvi2lEViBkMXybqeljHQlqpMEuMqqNnZNkJUpsdEgKdRXzp77Ra98K9NucbSdVgmQ2
94cE3jF9HlAOjufqJGZxJXe5i5NKdxVgytmSiiUXh7GBBU5QzqJz7Le2rJeUyiOszQ1iahf86p6p
AUg3+WGRHgIl03o9gYbb42YXSPV533PZUR1aLhQcLLphenzxa7fvZ2O3y1lgTYuxKJbFJwB4woSL
9NSFSMJsHR297uL8BarhFFe0c1Xak8+pxGYtnYF4/eZBbJV5VikiBIzjqxxIhL8UOwcS2W236kH6
fUnhRt0Cq8+QGvENiU/ITQHkbo+R1XGDQXrQn45ULts8FB5DhLYZzMZuWnN8O0Oly4ffXwR3gzAL
VrAi86+Zdl26gALIJovvvoabnh09sVoAvpOw4wt8zaA86vV6H1BvrI71zXZ2DwqGxvctjXgUvbFM
/wUiUYfPCGMV4pickFGppWpHWZ4WPIznN7wY862NKo7lT0YEa6woj0Fdn1/VNJ16UznL0IJoZ563
nGtEf57Cx8rMsIT43dxtR9nEF95uAyoPv2iTQqo1h7SOWi7G99EYyBHNB+xUKm9KRKe33dvwOC8Y
CoqCxyNQ8HNyOPJfu2oaSRgDqD24YO49dEcy2aIsEbcN9vq5CEAPWokzENGf65mxkTdMXIWbNzEC
Ci8i/45OQzYESkeRFnzeovWNGCvKfwIGXM30wNChFck77E8MwJngIE4WwGrS5a5RPmsnw+8TWFYJ
0fsq1SNaHXXPW735EhnnTYLT3Z8fQZWAKHF5Dnzg9BWIRE1WpJ8YBoJ9sk+3VEFLS0SMryWIAqiU
RxWAO7Gr7A1NK/OS9Ppor2Q3ha/IU3hQEr7ZjPpsIXmLqlpsohgpiTgLW+tsr/+5LIz8RQafmJaJ
F92rZ9Jii7QvXiP2c0St85+kGcSymRnCxeEQy/0qaznRdyo2oM5nlQIetVbmJ9DZn/nexipxiiGh
TXl/FuEQO53/yJsqlgInkQZXhO3swFs+CEZDF6LuSxguE+tbw0kkVAmuveOruG4cqIS/XrZ6SyFf
QaT+VvOdC6JESq6YmVR39lBLjT1+DGk5vJXYhgUMmDD2Lyx4samx4ETQ61a8xZl/M7T247VsP03e
8uMSfWK7u6jPPNN+EKBjmpkULMOzVYHmluqt8gzb/+p3EEtoqbuRL9tVJgfaLFcwa+tvJaBxer5U
ntIPiQXCmX1+uH1Q3LbFh+KHtrX1jMs8bKJN2CRzGN0zBUZ1T//EFSY3C7ESJ9x7c87uOkNiYi1I
Mw8hqL0Z+Mdso/798e/0mMxobbsCzG7vqmJh8+vM9tvSIBBfhHcHuutxqYD/6HSTN0gQYy8VOjEM
3TXMSjZR0Zbjo/2jp4sqyuyoCpxWD+lbPLtoDtOm4uU2RYJXpcZX2i6Se3lPBRdu1aABOH+FVvRx
kRh4TwjH/mmWbnb8fX00rjbfmpOhFfhBxXYuT+HFIyyfLMYkXptBnl/cR/Ik2n9K3QpGN1MTnL8+
U6pKCerBwFPVNDD4ZbORULBGVw/vxYfI+mmwQiKDIdIgL6H5pJBadNCRIIiBdxn/hmWpLZrcuRZG
/U/CvnVAwlNRkFUXemj6L4lmUajjI68iYDJBIWd5sloElEBMAV8Kk3xihJajoN/U5HH1JHvHPF9a
iyZlU+QiCtX1sYQv04O6xhe9NJgItNJJviofz3KW8WZINzoZARB6ZbmH5quA9+CTzMxKvCGj8Gql
H6ZTsesz66+efGRUdU2acsI8IqpDpxpT6HTEOum7XUFL2RWXPs+Rj+h+WBdZEir+wFzrZ+kPBrZc
NJXOXINB5KSgsU4chRia19Gru3Rx5t1uyqy+COkIulrDVE3ueg/QTbp1K2fHjzDe8QzHm/fTOkpG
b+5Tc6UCofKC4gdRq56BfCtImfHDsAvTpgHd+QYKcRE4k6T93h6thujlN0GAN8ArchMHs+AgLGfj
Ko5zyHAzaS92vTIxcKLxCvCp5VRu39jjJf3q9bGJ4VJnIs49Bd/KqBtXpWJ7g98cFKbETG/0A0QP
foxLpDQqrhnBJVCHVuI134KYDi8iXTQ67DG/UL1sj/F5v2Wc01ramxImbp+krlTa5lCVLUL6mHY6
GCTq+0OBuYJfE899nSz7mtCX9AT7fQEi9QSUWAIL+etP3dIZRr8lrQbFTZFEICt+y+y6yJjw3xru
qZuJFJHSxuaWjApekPRIgt/ZQ0rgbEo/aK5qzzy02cZXupqWVizw9U7O3CwTtnOROZ/5iNyuc1X1
NRnXKuV9LdHnzPyfYME3gH9IdHXmF3NdJ+ygTObrjme6cBv+b02RrNhf1KCGTUukXUeoOqsjsvly
0sene41OG9E6loxa8XVojWhvlBBRCRN22H+w1oJYzeWb1AxXQO6XRwHpOYbvadAv+aJMccpbgyus
xbVHccrvcbZRUkRetEbsIfSb6T+Ym5zm47D9CepzU1dY+rOsV8gLoCdtIK04qtGCuzkcKzwWoz4+
SXHnLZ+XLCoW/OegkFkjH0/Po+EV0PZflhTifY6xzwmR0oUv9J40g2cZEmk4esIU0cJrPAbpqm1q
rx5wjjptq3Vy3Wg7tVDOpp1A8vrC13XvZRtQdkSUFZ8jLXw4LR5mDWsy3atroMKiaa+e9ETiSTRL
T1PLYDapbggatvP6urBS1dhLe9UrTAE9X6OAGoYPz8m6JZFwUetDKAir/zPtCbvZdAaEM7aA20ZZ
u6pvrNtF/J+Qt9gu484+bt2FUbxM3r7pDb0HTmYP0MyOmZobnArQdHbkwnH5560HLDW9h7vo5ZyV
Mc/MX+1ndLA/MszPyGhnTKHNI1UPhZfaqU/eixjBLHOsqHuEIUDR5Y0kjjLYhk9/xeFOZEIBpCmx
hBd3A5UNhy/jAObNWJNT3w/7bQArCVaGsHUKRZDUInNMupMCPlmsihNMvxbTRlOTe2C3H/ld6h74
2uYuSD5T5unwlHeLBY5/EQUOnN0rkUtDBSwDg0VN1Z5WhipVXadIaNbV+nlK8sCW0sebv8RzLOTk
x6raNmf2Fe9WsuZIcg3z6oXkhv4aYK/9pfFl7yf/d76Vh7IOfdc94cuSL02+Qgs2v+YkFQEK6XMT
Q0U5GAfGkodQpj6YZn6VjWJNJ8SdB+gWTLlEZ1XJuHo1PssGL2RjEYfFTaL0c0+rg+MjyMASoDng
ak0ICCVi5qPRdHAEGbHWYKklYfqElnN2ndt9DolDlQz/kFEmKKoBEaHAbqe4xiHKDbmPky5yTGdq
jrwX7TJiKGq7fkMid0SwZP2Qvkm25mH+B9glynRbR8ItfzZvRlYetvB72mpOXDfAz2R7xal1Ih0A
TPl6OgmBwHiyeq0l0NCNekCDmTp3CZKMnEKvlCRFHYPPz+M/d724/q9Z7fi1H8N6mmABVqpPW8CE
GV2wPhgVnZR/J7a+WuesRFxLEkN4gBF16J2WXD4cXJFfwe785+4PotBxH68klaXeESVSKT8fxZkS
6eY1s8qcQ5NFH3Dfyy+mqJgtVJsFPggfVd4HPDmK+5gEEkom5+o332o7KxVdJhUXDb2Jj61Itit4
BjNh14mCvudK7pY3/Xd47hRBqX1ThGT1sMj5/ZmZ02CtqUeUiOsETbV9fTdf6pfNL+KWrmZgAbum
k8gcapXbNvueXmuQaU083VWgD9nwjTk/GvZlMn2kx3ANog4hbKy0laaiInEUbNEdlfSIfL5LPC+U
YstAPaaadNlLpLSw8+UMgIJyEOr5OdJsS3b8N+OsueYTVE7+qcUe5gNsQmi0m6pkgD5Jfd373hCw
ZF301xWFbqYHHSE987C+LQ8bZOlFcwwW2iw6WuAAGUHqpqHDRL3HqACqOGVG5FtBQO4bSZ7P9BZP
JIKnclaWWVjCuzgF6IC1epi+0sGvGC6EaBYUDYziPFGzLVaHMeR2YUic/0sYqfSUGEI6B8X1LZSs
vzcjIs2GQI3oqqAyKO/cLFG4TOzluTkIaDmBbS9Doujocbj6SlV6X0RqrBzuasoTlly5NY0tbkTt
+hOL79ChdoRTkHCtTSHrptFAoRdBLHtsieSNeBfuw5O3QecTOPWzMQEv6KdKW3ihLyC4b+JsgZHc
H9FEVyAUsYwjYjR2Q32OSHACVEQUsWq5x1lC2AraSFDOQrcY5BlcU364XeuTw1ZMQ0MioCi4zv1Q
AnCvlAD9YMppDKoC/MJLgxeb1HZ398EVTAqVXpNG7naIt1rCEEzUQP83Qoex4IfGItMPfUtGa9Lb
PYBAHJFtSsMLGAByoLSn0DOi1hDmPGVNRhHBRrKB7B74q4CppoJQDShokPZdFOh8Oqnh52yOXlEV
m/QgTyomvI+O4Oib6EEmlW8aW39HhVwCTn8n9WhrMZF7Xu02A/0izEEfslCSqIhyuEvXXchn2SOJ
8k/H9ZShd1Wi7LvmWszq91wTbHf/Dt+6DqJapt3M4yS/y1i1eOLBEi4tone0deEvondZ3ZYkbq3H
mrMaUrQ3tGuu7PCZNNMCEXQ+X3qH+4bCfCbJT3ehugb4LwASriKZUnhf3qKNwOnuXrWTaMZqh3gZ
pnmhuRJKagvkKvfB8YE6Ms9pDz5G5abEbwSgIFy+GX18JThtGseUDxUCaCOcyUzBHJjC6EA26zfN
cp8KqF+v5Wpm52t5iYlEBYg7hBrFtiYx03+/QE8K6sT29/tM91VdNZHbueL1q2PxM3p2ooxN2EZJ
e4TjEEySFLt+WtuQd9N8CVsvl9LfULqcFdqm8wsqZeD4nHP3xLjZLKVi262Rt6FPbOYootI57KUS
eENQW/m44Tifa1ZfXlIFosYvTfOsQ+oa2M0JMwlBjcm4EaZFbZ0axq/31J47oogEZ1Yp8bOzQRXR
glTCkJ0qHkhXzGNrdgQ3Sd8K3dDud0G6fKxCsBOGRWZ//alra3EqDlGdk/C35Sr++t0Ounk1D6xm
KmKyuwtafoTarRq0CnBWtmjctn3gKtYsGDXR3K/ib7lfrfV5wnN2Vky0aBEPi8NpHdsbuZofhLCn
uj1Zdl2HrWgoHmGm7pbMddvXh2z8W8s6NPyFn/9aiSeDRSdNwr35PcLu2x9CJDG+/CBcov4fu2wf
wWes2dJie1tf6AyG5B2y4rbcFDT2qIuiIy5uWZ/cwZwcncN8hskOBU9chAbcEdQB4Bs79XMTgFUL
2IwU0IKRP5XMkfIH12Syn4Kus+2nf+T2TLN2vqsv36eP6pxn3mYK6pEwwJWb7cp2Tg5LzvPYirnY
XLbgIuzrWM50ckszhjLdNF/KEiurpeRRdTEHRcTuhpf7WY9rOAOI1czuzB9jKPUPEzYnrv/Wbwc1
/4uaymr3vzq5cgBnMq6gjmKG/6PMnyrneE0km0S4hUt6k1m/nD0zjILujSBKFTNR0OYOaBE2rBvo
qR7vVHkt8eKyZ36Y7GaF0zTEmWkAWQw0+/ORm9FVMSif0MTzz5Soh9PBT8eTCI4uRucGd61zM0Hw
JPz4b3PTKC3BLjhu6bGmviPLCz+AMOzG8+4FtSYpDB1T6n0SLIahXO4HhPe8xrRkBTSc+rINboyk
TX/aFy8XiqobuZ0VsNCeTOZHqNinWVsFQSsRDt6muBfAeoBp4eSmyRwVjl8YJwzz4mzC0QTrt30C
iR6yM99cKo45ZCFCdtEKWUDWyt2xZoSUsJUz2c6mTtLN0UIrmV1tMsaaNq3X4L1VYMyya6jbrO4a
DGuImyzmQx3S9UPExg18IDqv4mKE+3ZusJ+nJiUW0t2s3Sj5LuaGk7kmo8MoOhffXCGsQaYtBBN7
nqGrpokHbRpEUf9ZaKcyxKBmAV6N+xSq+D1VmmDf6jdS/m4gkl7gdi+3ia2on16a9LzqD1mbCIZX
+iwO48GCwnQCWzHo5pi0YTVeVfNzZNdDUmj/UZOPWp5zNCpaaW5oakV8iog93bs3nPtu3w0SPnYk
gqeQiJ/YP9hTikWhkMlANZcVuuWfX2WxKYwmx7NkT8JMaAeB8eGZenC3IvmfTEbI9K/u+slDEGU8
Awd/QhlmuRLPz8PD8mjDcH9wz42JCflgeQ4ChBSdfq2I5PwDKCSsaJOWa2XZMaxoJ6tvI3Ul6g8V
XpZvgBXek/MRHHUrNCijAYyYCQoEXU07NfAOF13TZz3c09SRv01mbnH6e0ugHINkh+v7n5hLoGSk
0VkwXk8vX94jFu3IJ+nsOxaq6FNPTYEF67/JWtvHHz9TFzXRnXzchI9M7oA+sRPToJ6cFM3+Hc+F
KwgenArYEWmf2BDzJSY6I9ViLHl2lUQ7IRJqhprdNTiIRTf1WNIxzAqQn3yH2DZaJOvavFHxa9Ni
+28Ot/cY8SEvO48SQnhxJ2OQktp99aMp2gEcOUnMW4o/K2X5bUFVCH6G8ULwD6+35YGuzPA6IuKp
nXtWOQ7kyeql6WShztTlMJk5uYNf2M5iqSZj8phY1lmXp/Xof82ONoA6Ivr2TcrtHi+BFtgHOJvt
ah6SvZa8G3L9uVlyiKV2loVXuJ+anIX0XUcQh2QpBJ0+YogxHM1d97w9tRU1Pw1bimPJ1uVZWUQJ
RjzliRFsv5ctex/+l0GxMH3QzW+UPaml/wf0pRuUgIh6UZmmKKu9QIaOrtlzek2xxR87XAMm2DrM
pZLnC2dwshFltbHkUetzSVS0LZt4zvxtb2DPAN47uZPa4F+Q8EQ+TC/RfQ5LqCjoObVnZ72rt7PQ
2j0vAaI7tCaCCe37EAjxxpgBlVbNOoO9iwVDBoZaRnjithsx9KiX9T42jOVoRMlLTta0FSUYdFIC
yuF9a3g+xTCIH2JmNLRRAkf+aM8MC2WkxnS97V3QVmTldBk9/TBE+Eff7kTjekvBgOmS+sBdpNnc
OQNsJFwN92LKl5wwZGb34grxyZm5jPN0n8Nbl+RNP4UQNPfwh9tcwZRzKRgGT8CV7ENYiG0oIja7
OtbVCxlcsB5/StMMa2+KJojPuvH8BHFice6r93tzCYcXKFGi4Sy8sFS4asu2VLVRjnYv5Y2dT1w8
eTYuH32CfALndNPj1u7l7v+RVAlHS3delg9P2nm8LdLd6VonFi36GQ0O/dXtDjfGAS2tXUNx0AfC
mvZBgRBKfv9+zST7l8cvhr78UUKC3SSuZoVHZPbTCqoQacA7B9U7sK4FTlikq/QcktPAhK6d+MDI
qOOKoxseF+guXlCw4F44n6MbBHy7cNWK1uY5qBvdLRBg1qvO8qVMT0vjFjZoLIOF8JsLi6LSOLKS
ftZk7mq4lYearmDAXuQvkEgAc+zgc8dp3krmwZv3UAlWXvQz1eitovDtQU5BaSCoCAKg3TVl/Tps
K9LhuDG/eG3Jjbn0e5V9KjYm5QbkRg4N7Np8GnqOU5TenOumr2tcfihyU0uH7guaT0PmGniKI3b9
hzeI3H+elPqvf7hHmB2qQTsZv0OS4hth1TrsfLOVdvJYlN2S1nNFK/c38yovVUqDvMUibNPVURSI
8PKDx2sZMwI0Actvi3zlguxHhNg3myHJjtpSs29RDdWflYidbQ9cu412OFas1KXTwwZpQEuV0kWx
e0eZQ6T0DDgUvTDCsGnut04gZgnTeQN0Hxb4nlAHLy9ueT6R6mxPOWNx7H3XVScOkU+cOTeDZfUe
MaVswDXXV85Us7bRL/pa3BLurCYz5Ww+k88as30ZtYfAiK+ajU+dCsFLwN+ykeAZFZqn8PiGPGEX
5HH0bZPFboUtmOFKCdFlXTKAd6i0Cj8mFm6giOjMNVOg3htXVj2PHc5buYqp5vUBIso2kcaoTr7v
xZhe+9SxXau1ZdzTAe/IAS3nQui6OGeyCHhQKfq2gagEQvJmkAPMDseZsJRIp+eaWsMKqW5QKDgH
u3pSrKAE+rCXkt8yJy5b9GdE+SXKjfC4miC7/RnhrdnKphmjYS3R1VWfukugyz5cUy5nYBNg3S7j
T7y/SCTl7l4M3E0/2SqHMZQplLcG5SdM+II5aDpt2BKmdMiWN9ggjvUsfszVsi5RWn+Hfhn58Brd
I4euJ8LBtaNP2xP3S+KB4GgnnqGxmzacqeKeLPqMz0N5w9WBiMEzpOayZWRwzRmxFPvgRloGi3P4
r7YCNGg4ifZSvhChgkdS0wKxZsMP0OUtlJRy/3LY9YMCNu7xeEnsGyooZo+hPYS0ZPRrGgkCNC2Y
0LpJkOmI2Z3w9WElJCe72rZee6f7gNo6/5NNZ2Gqj+yGAE5hOovwjBxsbyarY+5gSpmtyQofIjjO
8hrIkK3IqNPFAhZkDBlxCFsRbfeP3HOSD5EEU2qr3WOfkLks6gg7J38YVvPZxkvOTW9K4f0WXQy6
mIm+zdigNAhYODaqgZkabvu+vbUQWUhS8LQMppFaxwDzjCqmUbjd2Ay+rnIE1UxuuKCkK534FEcf
ELmhiCi1kc6EHlV7ozPHERBAiLiy0PT/3MkpVBZEmAxX+4r4ukmNR2U99yFlox4G6b3PxYhxMBPd
mbA7EFqAKkNygvllpSbMsau0oSSilDJwhOkd6z5hnAhseadDGFgwpFRu0knPFQ9AGvq92yHNmj6q
O2FiUe3OHBlDcDb4KQBkxNhisXh3QLgzdmwh29/vblC/s7cWE/lJN+S483z8lwOkN0CikGdhK3qk
lfPvE0YxsP2IFPhPKCt0Tzfqnzl4cXERYuNSuygx94IQ995pwXiCc1cp/6oqsrwarwiYpxbSSGka
wFbdo+QvKSIcpCMFb9ANG10/yvln2tz7K2gnBEs3T6wLOsvatJ9IcDk59s/MmRjE+GcDCJD8iqqZ
CHuYWcw+fBmn+JKEvCBlxSaouzAcYZZla5TT48hagejoY6aALreB3NZTzmIQayEqe7fCrb5bf5OP
HxI7c+ESSx0eeRzrC6bHGWQ4BSwTzDS2dSKgplY2vSMsDVwkJzJHUkh7Q9cXdp/Jg73sTBU/cUvW
i47LEW01CHRJe6zPylCDZS/LzD8pPbxgEQznPHCfGPyNQprORqd1xgD0VfzAPXGr7IvmkIBsRfsH
k+bJDyLTwHvz0UzmOkQ/mV11AkheqrzVvA7A2jjZ+W8kEcj6cNHvqCagatkDs5oExUneYfjYM42J
xwrcz0r6x67KG8ejEsFx63kd4FE7SOURiurlb9xYizuwmISbkxLus1ipxgICei85YT0HLGqAOpVN
Wzg44ABmc4zRA3y89MbWNQ8X4lM2u7UlTu4eJhHPc1GhafqSn5BMQko3ScVRS+Mskq+j7SRviSxY
210WRAoXcB2cvGTfVu9FRXeSqqBUI9lTdO/+XT0h/A7j6sS/WmiWLmKCmveVrrljP2K+xOgpqjQ+
s7O4hyVqqkzRCmFq51xTNy9XI+oQjUzTzrtMYGI87KdZ3vah+c0Se/aDSQigP5dgaQbHWmIEgWDy
+5YPc3k0+p0EmTSaO0+k2CUxyMsnfwK480YAmmn8rwHbMl+Piuy9tS/HvZOBnPXS31XCB/VXcsG9
6GwF/0X1f36H7WK3XlYzZ1oPd9v3gDengWOv79jVQ+5bP66ob78TCjRsdVjuXNVnVJTgwSLFSDy2
CjnlUYc4M6aTwCp8pwU2qOEEYBqJadNX5V1EQnjpD/TukCmayl+60ofupGaALvU866/hlBa0pjdo
3dx93ITwBYrtXk1/ayEqIXCUmRh7dsqksgjLmlh44fqhVqQnJds6otG2/3ieqLlJTiguqphBFz0C
T7YwTMkX8qy9udfUVc6ZeizhaukZfBgXGflcMuppg1gSViU3G4WUyvSnWQQPnOWQNZUPIIXKmN0V
fw1LrokDfACGJeXVZ8iBYwGkV+CiFxBiVVeNJekeDEds/v7Ax4eVPTjJgvSvbX4obkWN2vOP+zj5
pMoeNuLjZa7XFJ8UUdqFzRgDqcKaDnWY+ftlHJlCCCX96QNFPIy8FBNEcqePG8awF/nwF6+dZTxI
Ktm/AuGugQ7qGdzBWTgeUqd+5FcjuKxIY4mTbfnX4d83OW2dUIlVa/tBM3+9ZZcyDdYP7ls7fzAe
XMHvd7D6ECC4cJ26uTlrh1kJ/aMNzR4kcz5ybKmN2xkNMF3TYNt9eg/Hi3yyhjwv2GVt6ca3XLpp
2HcDzl5aCPNudmAxHJwQwGj2YrEYHT4T0zie8qUuFXOC1Dlr4LYks2nkXOnp4MQ05mFDSOQDPKgd
pXMSl4+qEUnDLtDdjFGHLq8LFrFHjxvvh0SfBVHoaBowiLFvwZn5LHMhzXN6u6jILiPtzWXZKvM0
G98pAI+9yvrVA6qXF2I3WBd63qp28VHE3OSlmCloFM8dBPlPL7DHtjFM4guVp0vzfgN4i1KlTgDv
QGmBrTrGKpHzC3DORUIRtyuRLKJgHbewb0x7Gj42V5iwTy6R4Og8xXkwfYqqp0vtHdeZ8XnBQ7xq
YgCnhnzhbNc/+bhFkC/kzNI9xO4vSi/II3rbtyqQGXFRCPQTfP3A4U9nBCc2X4ZOe4yZ6M+XWNO5
vV312nSS4irJoSqGqOr8j8DohfpMZGELuqAbtgkpHrlEaC/8j99pK/ujA1QZ/ryCtKQIbaV2UVzo
24u7c41yonRjuo+PiaTpPtvPz+HXKmndeB4HeDQVk24VRUOHLeY4+dS1cYez0/HigxAB4IyFnSEG
6tcVK8RltuF0h6zK7F+6yPjBVl7pDocdJwd8w9E35OrQyRFukro5ZL9t2UkNImYac3VvJpVnBHBm
l3Bqd+K6BuB+zSdOIUFtyMYYmVQwOvBSxkyNs0ms75opuMuoByOuuDzaCjhWnUReChEoU3NyBZCz
pQHQoadKB4WXDjc//2XB4h6gE5AVfWMTkyk/nn2fQnbua5enXaAZpUpNxkLLDkd6ff5ijL/msvyN
sqjDHJfQ8W+I1wy602Lk1/AWbCXMsdjok0G+qKLelGPYG783gFMiO0jDTjbgnu+mRGbDVg5HqTHp
kckIbVkTtF6CHP58pBsMl/i/xezuTPxLk/JcP31+x8dzRHGDM90jtxIng6RbTGYKuS7rSAcLT1U3
MoCcJsQWhBm/4HTcc6OqzX/23+hFEJ37OzuFmyWs6WAVUwpxCfu47HmfZrksVOGrWtR9t3fM9a2X
YUYzbWA82oWIcZT2kDKVAOdEznCAhz0Ir/3go4hXJMPwk4Bc4439OodB4xHb9vgzSrLBe0GxgyBT
ufaoGOvs/ghi/ZU84WUNrSPcmD0H03FoG671AGpBpFilpWGc9J5rCuB1r4FbMSt1ktPWTrN4n+nU
liUIGyNqeOxUb7XBiKoqCZicSqIkiDcVsur01wDIa4xvk5w0W6c2GEwd6iynYdwYFm9Upb7hO4GH
cI/SAFYKRNThS3AyRLpRNivONKhJFVmnIWK6vi/PqYZnlhG4xe2gHpTfDGUl8w+jHJ+13FKSCfi2
9mLE2ywVHoAKRgUhpFjO6YHHqZ8xrJB+vF2KheylvMQLi3lOxPWjlvOhoQWfaOWeHS9+iAS128bx
PFOTmHJWTU5jUaR6GEj7Wlaf3FWGxSNIjPlIhRSZyLCat3MTiqvcgwYcSmAAXXmuYHSuaBBWq2xv
KHvAvbpZ69UZ8bV2j5zT4G7l3GEjguVhjGoCTLjBcT26qruQGKcfP3w1A9q1/jN1P+WAmz5zS2y9
TFz4jFHcgvi2q7x035Tiod4QPzmdcAC0lBPvxAb/nEURhTpyxQo6wXOPx5RyYjD2+fZ/XgXvgP+L
RPNwQJ5RKfL4Tt/dL0oXsnYdrryw+XvBsApgr/T3J1Ays6F95ePCIDMrP5OdKNQAYdhjZv7YpBCm
h9TaKwO8Oh5nF5MuIswOHHomLgbgkHhgsOaYeylNjJw7+kInU/3hp/mHkeK4mRhjhWAZP2iv6x9U
ciycbgwE+lnhV/CZHOLCTedNQu+0F8SMWwXX235/Xltb9Y56klzvbykeW3moNLvearLBU/iiWL9m
5q2fQgo3wOzDOKrUloqmQRIB+y43zTIZZrwSYZ8IndMxhXHhULk8cxCIRWjdbm3P18haRT415cWv
Ct0dloPM7adwWVQNTRexRYyb6twX9YNn3nRShmwIO47Uj723NRU9mGzfHN3ZR7rL/YcgI/yJlteC
UlmwczszUYs8iYpjb6U82tTSGrMUHg8r+F2FLCebIJqcJKX2QjYt4l9KoUz1EwXPm/6L7Q2ugifa
2BpfyrlRvHhxaepqYsLIO7HxCJAGMntML67b30zCDItra8bP9F3io8WOTNIL/J+L2HbGzNztUKJc
sXV5IuSjVKIBooQdZfaArpXLRYMhg7JKr1D83a7R01PmHEbaFOhLUkWj+KkxepWXcTRaUxeVfxlB
6x20Vq0rBG7/0xYnviXT7745UVzeiYImH7pwuTyN5wJZETbCsxIXM7keSjB55yiVM65pqcXSPI3F
BWNRTN6aWCE5PoEqh6CT5l3PXeuWV1UVgD3sZSpHFDHeWD1O+PbAw42BFa/H4Vpz65242jiNku2o
410+/+nkfz7asCtfCIuQt/qCnAFQOk/hoix4ln3TbfiNJUQQz4hTx6PQtDG9di3ypUEh5vn/2LG5
/WViotLqrG8mREr7FX//6EM54kMsOGrmQAMHpy5aPsKTRJXINpPTHlOemWD0fhjk4jrFx0DbIFBT
nKDmJLGsvg9NvIRX6pwDZcIezTvqAniybK1vVQFy2xaU2R8Uo7C/mS3P2wKWQTDi4fHXUjp/BvHm
s7DUv5WU2yAYAnLka+f5m6ypN5yb2AVSAvRGtZVYXs/Oq07QYISgSKZRY5W4sPmjDEbhXw/p34aE
Q/+vZMb9r01VuqziD9qUdaaHCLvYxHbBkwZsraEBhDbOjXw1msGwsogAqH1SrkPOIXEWo1oRhV/J
Etv0WIo/zx0IKlHHyrmCVwZVnYvQGeEt7PVfhu3NfIY60AZxgZ4s1SMqoGTknUlpJaHbj3hd2USH
2fbcWGh9ME7u1VrqJq56PZaVSXNrCb73gKbaceB5uTgT+qj1Bx7ZhlqAcs91ZHUQpovqqIDE3bFY
66R4haF0aIxeiyEnAMinxivGv3UCC1MKpiibqpGCJO8NGj8MY0nlDd5gBYjRGXAGw3Zi3C6RtQn1
6HoZJzRh13zAgMnkyittvHRSsLhYzh/ouyJ7HTj83vccuDGAf0mUbdFhQd59MLFsfRTU1PLOZiyA
hIUwUprrVOnVDc7bHlzWl+fpJ94TyFkN/bJR+4s4532Q8wbxNJMacyZoPhFNlVauO91md+ZR1xOG
w0UEGWYsUxfybfcTpCBWuSrVENoMM51GD6D+3VQzVpw+earIEgp1JyA8PoGyWTWtdvrwNo1TZlhf
wT04PCJhftxqplrQC4lEynOSSx28doQvkV3TJBuyGjocd4vVnMOTvypy+mcrpoJLpAFKbQDCjp2o
4Ls1ZMKFHrN5VbPdLu9rY7kzlTXHDdqifxid2oPD4lkizzLwUECeQXYseRUrn7CUu9jRgQgmfwsM
/37/h1bogP3C2wRcgnPQ2kvtmLk7GrEcNZ06MPFUubJH7Omxzf+JppQs5K9T6YpBwQrRMIGsPuaH
xzs0swv38nx1iuTn+obNfQfUoDd5GALbY5NJhl1dCP76yhd+ZvgZBMMpoXwK4DEpCBccGn2miqse
YAohUczkPF9OAWvZhHVjTVmk48Mk9JDuj4s3fFbALh23lQpYSAQ9LG32QwSKB5d/ZubSZm9w+epg
dVkKRci/bGQgCkfKb5a0shaXaqWt1hpc10VnN0Z+67Wjigw9lLJdfdSPoNIUirkTgUvFg0JW2b9U
YOtTeKCAft0U7klPgRsJYWomPyhym7vEChhZtIYv5w1pABwd3CaHDxZMkD5WJQ59OTfe1vmOFBNJ
EImKnbZHX6WAlZyd3tcbMGdhf2zDittk7tCkS0Q7YIXZxuB4nNJdXT8PxJ7Gw9tvhphs5xsMb0hU
MfX2dFsiaW+6uxDJ5f2c8oSaZ8JQHQXyfi81JnNuK4QqEgHM+hHM4+fqhkRMIyK7mP2skwKhU6Hz
qFf+Q/B98/o3wfstf73W5E+bqdVJ9Lb0glzlQ/N+OcxugdAiAzqxigNOLhfRdiTc1wCd5a9/n7DA
SzhPCazU/dGt8iEWlgD8dggnhBftfW5T1KPFQlAzqgnhG2Zy7cnUZRU7QeehFTl3iLRcMJ+YSmtO
MeF50wjpqygspmeTW2ftUbRl23NatrrcUNvBEHZoFaqTU6Du54IBrhMQ+PTgjdbRklE3QlzQSouH
wZmCT2OWj+mRjGaMo/uYffRmAC23LHQbnwaknLRLNAwGh5purGyRyPsQFJHrS7x5MYM9kl5fy8ec
SEidZk7ryywjqzGSWDMk1GzPEqYgM/dkUcMCyq5Yd64ld2GhYalU/qNGn0Ksqo6XJeHKQueDlSh8
8fHDFp+OZUPl766s+2kvGEzDX9grCi/QV45saQYd9R3gl0vJLqOV+d4u0jzxG6f+NvFZ8kDS3Qvl
pCXYd5LvM7e5lfae7WxkigOOUjAx6HjT0mAvW1AorLJ9xlFWwZHaOeS4ByKNrKoqE2TMFybHA+td
Sz/qQn8NxFkdJ1HE5FNPdTRUAh78d+9K8KuuK9uKrxXwsgV2tsDvn1I6WF7w6BHg0LNnFav87p1S
j4ZyUrRTbairLtJLFtZgTkrnM9gWk6MViA9r81mKKWPRVUfo8zYh7LNhC5zqfDoO2k/tuBs7GZQX
p6wWDS4O+ZfKrafEg1rjCQSZgLacDfgMTt1PQN7J8Eiim0CMipQJPalwyI519HjyEpm/faGKIVCv
CHgDKLvIE8koRwFjiGANdbrTOQoDsz8SCyNjDhReKayMGl6FRVWpXIIvUR7mQp2fbH5oXI57LTQj
IEOW/InvHecINnQMdJG3eThA73S5jYaCdqA43C6WCJ5MpPWn+634s+AjuSyYrMcAS2ZHyrt2AMKF
U/38R5eeDjHE/cg7UP6do7dnMoaEGZl11S7HBRazOd4a6uT7tKXvtPcL2hvbRg52CyQSkjvOO6nH
fvR0PWLS2S+pfZHjySYxObFBeI7cOcPiVVpKd7hRdQaQb3RtIoVb3MBdl/pSUHOxi8jVRrM676Yy
SlWdaHvqOp1n06YTdBQxMdLGDcjQO+4G/UzG1fPIoBolzzIv2YiVVtiJdejnBGiCF38w2ZUqa2eu
Tgk0Tgc7U7PTDkCYgw5r1F4SiyIGbSRD0XZo1+nw9WRrgKsGF3bH7I/1Dho+0Pdo4KKQ/6Ie2zoD
bntSKsB0OQ3sqAOZocnB/LobH52RC4M9rKr1K1VuQ0s1Xg+qmmC/S7VXQnhSVLfHGbizXWwaJEWp
IF4K6ZpOiuFBPTmvaMiE2rvQqbBoDgjWTQ2nO7s2XrbfbNAtCrP44PezdvGVMA1Ci99IS1/wlQsd
O+ME4TFwbJLNiHAZRmFKxzc4cqmPQrduO8qKbLi/MPzK0uhezOhmaU8lQ3cFeKQALDUd7FsOCVGE
vBTZap503BwXMWrUsbjuLm5T+jtUwcP4nDGXBifsZSvVVjfMdfj3aNZ5ZrAwthG9H0kHzmVlDPiu
oEvZ2HWgPsIN9c7nFIvPesUVK7WKUB7KCCDpmraQAEaZtaDMWry5xJvcNLJzs3VwDxiby7FvwhlX
uEdf/NAVYV5VahNyf3INHx/5EKHNNZ03WMpx/EY5VS+GUcNBRnFTeh5kqFevwp63pMIe+Tv9tVWI
iotrI5HeD932AthilbNbaKtytPJN+J82v1rceJn2qPDxumYlnsSLW5ZxoQ8uMnx2zzAIYoVZ4Dy3
QtM90U7wme5Bfn3k7ZCfXp8iWbYDkH71Cnu4n7Ycln9lo0fa1UAhfBegI1VfNuO5L85fxclm/DE8
riqMsahPhs8bB6RK+qM2IGfnODFjhBmsEjthliQjeQLliNu2krUUyPYE6nLbJlrHiwZChBBxZusj
zK9cBXJSojLInd1SSgaZLyfOTeFNcS5ydvc9LvS30Id2nHfEA6JFFkukWM2Gi488PVdPT5OCJpMM
3FQx2n70OEoLn1g5g1TfzHh/6Mw2aVecMk/MlzX8ZMkNaXZBim7L8oYMObRaN4DuvR9Zx64JdILR
YS+MQgQ0wwXJzZw3v4L8ZqxFl6/Z7uDVsQ1bAsDAvsc2BeLeU/nR2NIrrR8akJmUxR/9OZichd5v
GW8durS33FZyIZYeO7tUl3kH8v0V5kGD5xUJqfCuV7J2nkqdYurGPcwDQS1pD+Zr2JnkqIfaoJSW
Gy1L2CPhTlvrlZDZynErVb24qrC9L46yFq9moLMmqV+qHWe7WADYgatIkPE7qRF6ZyS+k8PqlpvH
vaRXNxDg+GOe2uHl69FLhdiNwoWfo7To98D4Jx7BSygBcvcvuOL/y1qhv1veOyScM/Srle/jS8vz
wjqVpa0CyY6CgSP9/UR4VTrDjTjvLSjDtmF5i/RaLtk9TFmZGPT4Ia1AvsdokY/pW3IMCWVsu212
T6g2yWrUauPWzNrrWC55JqvIUJy8/EZ+JuOIRP1N3rxv3JiWi+1/OjtMT5745KDARgHeHzmUfJ4C
0MP/2QkueJtVYFejCvJrdxX5ATEK1NIRviMKQJNvYokioOexN5a+XGlkcAxjHkcgn8n7jn7G0NIJ
Z1Yl9Vk9U9GFhKog3zpNvVFZhZbF/GL3jSd1xDmJWngCmZiL11KF5aPUFI2w0rBkZusiZ3Jf8yTa
y/0R2VyqI+dTbJ76XmeX1l+LW8dWZwEvpMkH6MrV9Aj8H6f6IkHN/6hOk/0RAmULtcltOVDL1bhi
Qn1XO9RBZXyESiC7L5WH0T+E3n28e8EGHZkbdnGrz3RPMm7VuvofdsXxV/GyqqUDcLaw/Wj/pwr+
YiRVaFoCeEPN0BpM6MYOaIdCh9Ksg1QZQH7VD09+amOD8dJgWq+ZlWsl7/i7nVZuTYimSMpqHbHN
Mb1VPKH6dIP+c5iF66DJc+W/SdNkyKbS+SzmuLsyPyp66QVkJ0lTjY95IFo1pAKub9l9BOjMvXow
Qawfae3iXfbR4YX18O19cDHT50k+uVdkt95bxRD425GR2B0U6MBBFCxSOOaVjvZMGH5zXg13AQwC
T+W0tnJ3ZbrQNWYGTzmctjC/pViHe7I27TeaWDkPsz/BWkwC90vSUce7aP9oN5QnSRZZGaGe4p2h
LLsb02GpcQ1I2PbS1BIz9I2/pLqLnGL4r84Z6JMm5/wd05fDVxDR1jTnHwSXzq8TfV4Rt//lIAok
7NzhbJ1kxoQDNatU/Gmfz0sIYrVQ1e/RIiqPDDeY90Ug3x0sHeABoXtUO44lSdUWeHL5MQ6cz/P/
XIe46jX/YFXu42funHufdbaO25l5gHE+eSi+TWO+0HHIg1NroGzRXt3jFYo1szvtp8Y1ah2nvQi1
Pkx6njhRC2myfvfuLrrUwjsXcgO5pIMCjag7dV37r88o3wM3G/EHtDQn25Z/XSSloBV8W16jTjl0
twFuFj0Ly6YUaInR2RKEk7BXTQhZPQ55M3WYe5JRurJxS07+zLohdlrj8OLojLE3RAP34mJBExla
/t4L/Ob9kFgciYAeUhJd3jMhoJLQllWZJmHZ8xVRGTkZw7qJ1v2EiJiH6yXTi8n84IMG4dS9/TLs
b4oystKqLGcZkQ6ss1y79tcXDXZvBK34DTYna6TM6AJYJNsKD2jUXZH4c/8HL4VAOJBxgczN6wTy
PueCAq8WbW87gN2eUbSUotqKFfUWGJ0abielfQp+b6jWgH4m7pQG6YiRC9Sv2Keit1JJsv26dOYc
MHnQXtoQ4Gf60XfcKRIWzIUgBX2P82kzgLVl8ukxz4LMavAJDdQtZKwY2KexvzaZcTe7mXdryxyT
2Avo3g7I74Kzleel54FmW5jaNVd0OEboBOcEXpI+R5li1fDBk7Wur2gQdRoRhiMpY6EA2Qqd0B4J
HvJHiGqJCe0itel2HogVSJvsbzNVoh/YvMNQZKrmnZLraoewOzlOfAZ7IomogXoLMf79z9r3wS1i
ywvx37RU+1kv1UBQVrkiTfqjDi63fj/b7t2eVJkAtxhO2PS+u62qaObmwVk31WCQCIRodefBAQHC
2M+ze6lJgfP7CJaB0W8SxxU6ekMXcl6cQG4XSkikBKrCSc9lfIiy8imXqZn+kL1AjyHNUQ1BVzAw
g1t0tQucYBUGeCEQG541mBOuxyHTPs672eSAISEIPqVWeBM8Cz90n8D+ykt49s70rh/35BvxQVYs
OMybTwYyyEZgr6Vnl24D2NSoMGx0U3eFm/s+vlBV+1ZpSXobMZpX/Xia+56lbo0vhldyhU5vtWEc
G9vhd9doHNsF79zRMM+1TlcDJ0VMwr7j9W9jO5Fmtt7kqaH6TICOu7WlL8j+SFvKNOHG9f7lQGrH
B0nd+fAPs6szK+RTZSobjgnWAXatigqndGD4EBJHwtf3RwSiwX6o/sO/9GzQJblfReOaSReyUWqB
H7G/IxidEYNGDEceUJYo74zoYYLLdAtwUPARsErnIOt8usPVBOPXxYTDtP0tQfG9fyPsmng3Zaoj
a+LwgtKiWtxQgLg8OLTFh3W9fh0WqQ6Gz8HF3hyFumrGQ/oYPGn6O8ynG935kSAo14gS5YbpDbUk
0UFuMUDwwejl0RBDfl/5v6xqVvpD7sQSApNzKTIqgtVyizFPTF3bACCVQc4dBw7k1sRUJEV6aOW5
3UruMaR2VYnAOwZ+at0yIH2/yE8/4WOCD/kNTKuqIS7IN3+YWCjxBauu0SSO9BDPr/Ph+xnYQuau
ehX3W8z2JSRmGZIwjPujMJrwaFV1rFPdaKIwWnUp45dffApLMMfrVqt1IAghFB/c89dzuiNWWix5
UzlHdpbCDeYeoUiRCOwLgVz8pFxoOvuWii0nx3li8REKGOyn2toYyrjYVjo6R3XTSDSyxDiK2EbU
bzVleujTPTCVcjRbml2wv7rEmCx7FlEZfimZlJ5cPxut3Q+cDzScf9XxwmyOtMjKYGKuyc9TF3Ny
+v31mXcpMF95I9EaVGg+T9URpKw1i3+zccsVZVpXCssCdmPKBqRT4aumpDOszeIYbHuhDyFz4Eh7
KCuPOF1Rg48VaunFlDS+gc0LekLm3emRMWdC1exHDJ5jUkwExipIuC2RDkS8DQHDin2TdfGiv6km
/1QuW3hk6+BISZW6m7q2PkA+2gQbwW/cFgnSd5jwJtV53FGffS0xBOjOE8vp+degdolvdsFcGBlu
y4p04kAjZrUGcNxZY33A5uiVAOz5a1uPMYf5326jPNCLlxzVDLmtL+Hug9XN2DPXvsBGrdCpOpsl
Gb73Go7Yf+Z2iEXj1VzLt2ULqtdwYN9jTRJDfG/hR69SL7ilLwcBfo0LFvvAa5FeO7hIgom2AQt3
EKFlJPd//1XJfgJHhPVGiRGtzAnr+38nt63Am2LmDphjWK1+el7b0xorqIk6aptZT0sxWEiF0pC6
w2CjYZLo47xsYbsnchlfKST4Asm4b5neX99uJ4akTpMlOwYPQzUMVuFx8DWKPeZMkO4MLElLiViR
JEH2bdfm5pkmUJLrGy3/FFCGznLMZpZtXP9u8WY4UXXMenA5FX3oknhJy4LMdntkWE0Dp+jQ6+5a
wS+qndg+zJ7rtnG/pCGMg3pMZ5q2PGOJUkS3OgUtwJ1EqBGmSPrAmcBIeFFjCCEvpp1VKzkFBddJ
4nPAi/Sp2ATH2F/AFSCcJG6Y8IvVrCnuNzToJKr/hGrpZZQMqCrk4rVUz7p9FePgL5A27Ut0Fm3g
59Ms0aSFlNqZGu9YFe5OSgsPl+5JZ3cjmvSB22WaX6XMWxnfuTs/pxAymZpYlsESbXlI9ni1hOKX
WWYebtEDpkCGHqqF5kMUXn9pNtiAkXg1dyF8q1SROBYmiJ9e9vuu+s3aTWFp11R3jkSgBvH3a0iG
KXCrus1t2b4osXvv/SKuDWyhbx0OONL2ejqaYzjcsAzAope8tRzxAeYCLWQIgFHnWYSVFPFE5Dc9
bEUvmKeHP+X9sjX9uYbOMRzvv9hV/niWftNCRlOe9HkwrEPr911US1HBKqJDl2YDWYFRq88eGUEz
JSWA7J7WxNuV7wXg1eNatufHHZ08zMnEmuMXLIOL+k2p7ssUwafcI6FpEVGx1RyNHde+zJa077V1
WE84BKgA+ws3UpOVD8zDtB1+tj4SmqZyObYyXd9l2SWfC0YbrhlB42PKHymfRV3IGHwZuDTG/Qn5
bf8qyhxPA2TyoZ3kMTnTb3OSRAIo2BGgjkL6RsBKOKzXT60p6/WrCbQkUenIqHmXti2ASvQrPpt5
04Sjmocqco0njdF6FxGK7UsSORXplv+GXCIhSDVBRuLA0N+ZulOpBOYgG8DSvxiZ7jTLYEhNzRMO
8/w9BVqXlHI8Ktepzep+aYOkc/l94xDKzeALRNneQW4sUO8mFus2x/d/HKAlUPprDukAGj5q11rz
yubYn13QVf5+iW0Sb4A6yDa7oIyGlRmN1Zl7gZNPhbhTfqvIWtw/6v2SfZqu1W5Q8zjHtcBKU8TD
Ocp8wSl9HkZeQSkwNObw3X4HDbqp1v4wJCuSFmVgOjratmn2ambPVD6a0IeVsN24+ANZqvZ7N23P
AQlJYwbE4cl269bwh73jxvBgh2SwIreRm/H8cyRXqdFoR5HrB0ZPn370KcHfZPg3xNgRxanOZZLJ
e7HZnFEhf98CKH48FQ29fyHJm9IFTyp2TQerrJyiUMs4P7ribe5bLbLtHiWI33Q9vUb8T8AVoRzO
c4+EPnzMmxUOwXqcJgCq8PD1ZVZkzgrf+Q5Z5E1enecsvhHj8d+J+Fd5CQFrB5qd6c98NABrl0Jt
yAdPqhkkD0rH/p6N07rimYPkbl+4DdjICRPeSw/YKlC2h1QMnCVzhFr4gVurXhZ5CsfLnLBWWSgV
kZuo4+XBO2aIl1tophBS2er1Gund8ndutjTMyXgrvfSvIVgqiPQZHpTmypDajm/hvdeiasuwFkCz
2Vk3nUX6LcTTqqA6+PZbjIyOZ5/fmuaYdGduaq84qHMIx3V2QPrixRKfD3NfIK89zN+KfnRUMPQp
+tsN9l46/l83kqRSJ/m8C6Wu5xG+6csAuKNxLjvscMWt+UhsQ3PRb047400WNh54lTK0Mzu6jIRa
RcaEGZRnpC5tuRqbSzxruPyLJCa6iRjCG22E9V6+NroWDq71yI0u3GITFISlG0Fr/tEAhvBpEw2J
oc5848vF9aStVXwH1GV8F7o+FVo99zuwcFpBxasdvnqN1meE/hp3U1E6LMkA+J/ejfO4VQujKkdA
bedh5SXK04kOJtgB2NlTWB9hvNyV8RzcDfZCsHYEhDEI8KnFYzFsVnaLOg0+ZWwcIR+leb+2tt6k
630SZlsyjWtcj/iKSWjiFpDYs/gDYRzrkv3Hf69cvJUsR1YXtRRQbk69OcJ1CXbAWpyKi8KzchMm
CkjdIZcl5D24a/9ANR4d7ofrI9X2YT9n2Z0BOKUW9DxH8IQiYccgWHmflEl6vV3P6rcAxwLC2gm7
gh/+rXDL4b6uUIAM3KA7/yLeSWLd8tlQGLkxGQj6i8sxf+KRqPnKj3mLZM+zi1UwbHu5pavkmbZk
Sl4K1web5pAfEVywLN72BMyzZ5JMqLqsnvXRudnAm/vSANYFPUZqa7jpvAlVeTFUPWCY8rABOmXH
otj+C1wB7mLawHWHkSPvWEPCpJkUrewIC18YLXkHzQtU6SWGwgFLEOOygeq4uQB3Zkyr2C3vKCe5
ugtN95O1cqJliiDJrbj/pIz1XEvBAUdZbXoH8l1gNsmHl6MR8raCL1snxTYy0RMxT/1YP/Lkz9HE
3aUn5V5vaMWzeQFnCn4O6lZK1Lb7Xxh9wtJfxucMh9a5i4OJNGpQ4kQ+zJ5hnATvDGXouaWR1zEG
jKG5THhlr75LO18DjJS30aLGAPOHwUmsF7eXHsvC+yC7VJmNJ9b5n0Tkg9pxUMysfjddOEozZKcQ
0tAccW53DEcPI0wqeRd4gmvUcR24Su8CWIEA1nz+P/PucSN5jpWa0fFkqksity7Jqg+IfBsRta5p
TuKTbAmT2GXMdvcRxGZvgl8YaDerZy39+ncSbQ0go2lxq6arr/VsVW5RA23entuXIz2l56s/KEQ8
XbalPQRfTPp3/U8kxouBpWWvZ9Be47dsiNR1XdEYI6a8Tz3rJzzUClLZOCiCSGIwwwYeq4Ry4MaK
XXKsJ7w7cWPgJ0PQmciUzXNWEe53OvrhxiDVcczvBeRwEZnSXvEqN1osw3gifJoTCN9fsrpKuPl5
dTG3ETUSCf5Fr9OxJp83p4ehlUOkOsTrbl3XrDTBsX5aFeGMlGbFDBVI0G2chMO4T55PgxdTUkjJ
cUzuh9Vte0c56sD3jfHkj7Ijk7U3fqxKaigiqKPV9ZzSZ9BpaUCjeKUmql+AzMHCazpOhtPhrs4Q
fR5db4LSm4BjSCoznQKuRrX9eyQo0MixJpQzA/ceNyhXpLfMTBc0BoVhhSX5E8PEfXBCJlbQDgfa
oKV8/C8WytAP34m7yOcf1qNIhRUs0VGPOL7+kh9LX3YWy1difQPz6Q05UgX6ium5+XpshghVSt6b
K+UzBcRNU7YbQQPo16eJ+L653f8vYGIJQCci9QmwNOO3IRvpLC6dQCDjpN/Z5qBBGoBNECmuUt6x
AxXpJpTXu1o2Wz4b9agUkgiwlpFKfuPqzyNfl++RmFgSFLCnDETDhPFhoioN384zToNnMD9Mb7sC
w9ua17HY+W5ZiV6rD3Y5JpoWP08RRREHYtDUOaoRecRhQndy3jgDxmUu/zqJox3GS7QWcz91dq59
bU5VThCcoarjP4gIz86WnTWCZ1XHMLy+Vgg8xWTBmyaJ4kxiUtXsjdcZm8i72xK/uFMN2XSn7yFl
ee9fvix/AotGGlKAsx8vu1vUKx1FS69txAFOX8mUWtvOKBUVH3PF5yuhv+3OQ32W33OLptZ7ijjL
sMj7M2oIMi+3crd/R13Daum/wGh0YsnWgRLZaEPkV8XUGqxTNjW9Vwo8GwAnEfcsxuqao9BLK6yu
ukYfTTNfwA2jlqbzqqOV9bebx7my5g5Lc0GuAMv1Om9jlMLJDCAiYxqiuqUdFTzhJLapn3+mAJwn
ekZpV2Pti/5XFnqIQoi9YRfUS0aS4u9fr/bJB8M3OAF7tpXXJJG4FnocpKF+V2Ft2U2sPwaX9r4D
AAaHhINdGM/DMdlAk+0O3Kviasu02NV6t8XLvwZeDMadsBEDwEVTrY0aDfxBgGiqJrDo6cy21Voo
+6DvYt8PJMeK/l+sq3NINxoBYtOdEKuSBJDWxDqqKDcdCKBgDyNLI/RD9CFYQxKyLLj8HI0r7734
OLS98u5tKGjPVG6OSWH3Ly6Xl5B+SI9tFTjpMqykzo4TuPL+0HcekVSIhnaa3WYQ9qkPYFE/tNUh
3qgfVJ0Lhm82m3FTdNzZQp5akDeCDTbrySgPGNUjAs4WOwjElf5WJ8KrVpyFxpTlV9L3K2thhFUd
mBJJk77/x61ViK85Aw2aekNHhW4dz4geC08pThvyYMsrGg4c8bJWixfJ9WK+IJNMwPrUgoKjbVw4
CF/eWo3Xcyy7t09OtlXT5Caac77Yo6AhP/iA7/a9qZnSsBnSOp140pmGsoPsgL9EwJIf76rB7seO
HNpeLnmY9qA2j26SlVklA4qIMx7Ay16HEhsptmEe4nYuE84xYLV4NpiN9mIHnUpjb993bfX0TESj
GHexIQxc1YwpA6yv6y1kLMXpkFQTPqeyRpcGmXhhGhG5sCPpegOHonTCzNkxja5pCOvO8ngJsY/W
I3vzb31BMHsP9cIFvmP0CH3nzbWuLZEWlt7X+04J+INOi6w+Ub2dqwy8oXfBzYjveLFsZVyOtdOT
N7j7/3lVO2tG/WVXPDF/UIC6hGhLRe9RedeR0ZZRQRLpfPPrXZFr2xdYxjId++C83bv7Q+ZrfBW9
662IHrWckHBqjg1WTQUe1G+ij5bFQONmMZnRAF1q9wHSgX4BTTgEcDZrftPhSI3MfGpCEIWAPz7M
/YO0Y5MbRj6/WTTVv2P2pZrJ5uY7uF7OBYLbT9mp+fQbP/D7lUpjWYFkTfZASve9h7Hy4Q83592a
4MmH4Khg2ich4FIWREfPOlwTGQ+2TOZpwpWOh/uhauxyaahsFNmNHLiMGhG0aWAAs2eEMTsu4i7z
AxRul/IkvqHhcZw3OFlok7ymApdW+qq+XYz+Mt8/mmz3caXMTpTCCoZ1wEW2J6861w01e5emFHN1
CJaNayUNL8a050rsFt4ksB3seXluMjnDWYpGnTw4g9eWW0lmHcD9dA7QUD9HJk7G+zzJ380dKDmZ
KIyMbISCxT3WucIJU/4KEnjATSVzzXfUGm9/Ph4tO/wJ/kjSdqp5IjTbOwggxpqOQeBxdt6e08WC
ow9haI5RgsU4BUoUR9qHWMBfgaGyDBfJZAybXYK7K7JwlI+ljstdANSgIFXxJrGUC0Izo/eyaGl7
XuJcAuTDBbzWerN5/fxqX3WhNVomLqbNyiiZ4lIO+6NlB8ANzeXrm/bKshuvDWnFV3YnwdvS/X/D
I8oeuHnt2X7u9oO8KiQrF23hCGwGMEr0Z43xuLF+MLSoV8Q12DKs+XkLT/iKuiEMHLyDeEt5OYUQ
g1l4bijl9C4zZywS9cw7cHNcXgS6h1aOVwyCoIXhU2M0vbaGO7fOi7zarZg/JUMBpcKgLnoOaGi5
t4JVPqf2wemDmZsP546DGh3uTKDlTyFizpKVyzWjY+bqddaDSGd2aYL2E47k61Co2N5JQWnZdyUH
9/HropmfWTIYZOIOJE+QFRWwGjpF3mz0fhEmwny/3+LZ72pX6OOpOefjJRLhhBpG7O/0JawdoLQD
dIeXom5M8tDywFKp7pjujFNmWPlVxDnhvJzYzWTftL/CDNlt9GpZkgxvz03QcKMoVHQBosWjTBn+
T/TxPePU/5oTmp5RDhsEo/zdtH9bvbeGtKTuQuPXByDq3K2OobRsLviYMBMtvp8/8E+/WDDwy3qJ
xz9SP1DK9QfSFQXs1qpJYwB8uZSwo1iqrF/LItrFyNJ+IEQAIGxMMZ2lQohxtDm7TUWJU2UKUC5x
nG+KX9PNGkFhZm4fLWAxoObe5kbhXCbXJKSPioU/suuvvKQPPFGJpdnSdcRynDajrMswQNt3AwAX
hqs2hMiWzR07V/HUYxkhr08lHiIAeXnKZ4EkL5S7fracTucIR0J24OSdyUfNC05t4zVr+o8wgQIA
fabP/W6MPGeiyhM1thni6qTbEKn5s+g+5ZN4Jq01ndvln3f8Qfcf7BGvpN9/mKxwgtUdB7gpFpwt
Ldj6NqMgMqG2uQyGSfd8PL78Gk/FqZy4UCgipLOaTx5XUYauLOYzguFRe5J/qKn8YzBU7PHu/ql6
CfSsdh7OVGZnWosbvNrqNFvvpg9bw1QGkNoAKeK2w7WbrlLsMe1XkKyRDbM6X4SOiq4eevvnMIqg
lwwxNgULpBUbPwfqme7tp6TsZwlCDuiBIusn91HNi0rdq7uvhkccKQKofaWi29ogg0K9Zf1DP/6X
7Rr2AAr8MBsm5C3onZCgdN65RLRGH2ljTA0YF3IG8wg8+I9p3f4SdBi/jqcq7IpTk9RiY6B+gRNv
U44HaMGIFjyx43KuA+Fb2+6tt/wROIAy/IBRzdIE9FdZnRv/zYCLBZVXBjddYd9ikeLZUgI/BbZS
77QdPEPBcJekjCxakW9dzOKF0yXQyHaeTDk0tmhOydnkq2lX+viUR472qBtGm6Pd8snXbFDYyf0t
wimYy/dqiXIJPXmRs6Zrg73LEnSfqkiAbWCggM/Y1Z6HBhZ4Oc/n+QiRvZetef4XHPnkwRPu0sn/
H94WJCmmqpo7UEXDn2lFiOUh/GMr8a0Noqcla5Fy9hr1NZpY6WwWc3qYi0m2L7Hx8PEVgOGuLHgL
cYfBlhd4sMpXincK9a3bmlDmC8MvDGtRQ5GV+rnJ7MGqr/q37g5d9LKbfZ0eIgqJG2k6ire5NE0J
cwvVajALSe74dXkba9a9vCWciGBWtt/u58HMgZpm8iv873KXwtQs64dN0xvzv6yXFtwYZWRJ+phE
DdW/OOSSbf0r1Q1cZw0YMxIweJbq3Q6NucpFrGaH2R/HVXj+xqOHvOgzlF0S85eSf3ljeTpmfrJu
kldVLv9W7ACZLgcpfgMYPfpZs6Gny2PCSL4ZP8kRis9nzIpS8N6MJ+6Sg8D29F16zGw+Byn5ys13
jWnYY7hinoo87RKeaTamaI8GhrLRFn8623b36HnJ0Osv7Y1G9fo7BSX8Fs+4iIaSefEHqTQyXd7V
fa+7DW1/BRyeWMXH9dmUd0Z/P5yCQedmgrEbhnelb8sHfYuCp7+6L4bApIl/Nmxe5FPsksWeBJ0g
vCLYrWgCyhBuTrWf+KWx3hEiaDStRMQnVuM2MEvEL2MFh3lZiBMsnf+PbQUR/BCmq+dItD05t1Q4
hAG7FSHaCqO6+XZel+odWNDrqieLrlJSLJ/jH8N+DF7eYJ8J3hFRWxqr1YzZPKYmxwH4hpz9qXdg
ldaI2hXM5UUYhCViNuxwkKRav5y+QoGDDJJY/UCNkmOxaFVQxzFKtPMr+WBgCHuK2E0kGxUjJMhm
GIQSATqpPaTIEACYjY/hqMcmL/cOJw2aLLIEfuuD4I3j+tAt2QUnaQYutF8Kslv/imGX2BPPUAam
NDsQljN3jAEhF8Uin5cMEtyKyFPChbESa3qk9e7jNU+I4V5sP36JyL6tiNsxz/1G/MMxwZJ5038x
7AeOpXCdknjPWm2hOW00zRBHt6i23D8knZXzRig8vyNEw5/WuVGWDvUJT3J50bv7pKJCCVRAaKX6
aADHppk7C46M/+3oAsLF/nLugC/o0aq/Kd9y8sZVw0yaPaAr8tJkRWA4jyR9nc7Vs1tKZ+zdzN5S
M7nlTavbe+cG2CHxJACR0JiCBKVgCFMc1gFxPHo68dV6VINTcUJesCPPWqMj25h0wVbdujFDqaE7
pS92f2iUsLKKIJGwtASqP/sNZHhXeBEB99K1bDcMjslH603Usyfu0DmRwD2bzNrwj08+fwHkn1Yj
pkgSyKpzSikDm0DNaoD3MYgmqpmpafFF0ewZnf2a6IxaBot/5LUAq7g+gFuUn5M0/NQDHws7byID
5r+h9/N9HqUOMG/YX8P3T5ZQp+xYrKKau1gsO0LAE146VCMw0vjUQr/zHBITYWjFdVm/j3iym8QD
PgH1YZAfEhIfPfzBz6iaoxIydUVFWXGOgOtiOZ8HsYOVDJGIOD6kXyDZHmJ966eZGPf5FaSvc7+K
qoOvNvvK5sTYcTuQrx/mT7Vzfb2aPbC/20vuTwhq/1/wN6h4RDKwaCBzL6sXw/RzvHRkoqhdhS75
CE3aF5rUn39aJxQ2JqGMSDvDGfZitPpeO0gfr566yk/CW6IqjhpmDk3eEaQgSCkdsV4Ky4eUpTID
BPm4ork6wRS3364NWyaT20p0HiiYXpw9cQ71Q/6UBfKxIlARBG8GNvQRAXElLoweHGw4jTb/+NCy
t77lkWc9ntcGWMqYrd8KPuJ7jvwYS/Cq0yjyhyQyXjUoCmh7cbsq5JpVBZPdRvB5phr8pZUYKrwj
votuJX1w3F7Hi74MbrU1H+YelKBhMquT6dE1fFCjjnf/XThDhWYTsZIG5qgKnRoVljoy1ukg7NwN
zxhWok9lKr877plF1SrGqwgLJraHxJtdq10DwVgOZ1ItXC2uMvEaSuR3i6BH4tY9anaqgCaQ2ZoI
JUnVSZYP6WTbaFf3doYnVqRVZRIOxGFet0E9g61W9mtXYzjI453EBcYESnOEDCp9ia9ZHyrfrjxl
1RIylEPIUWcoWVHVl0VxpzRUzPkx7dwvYuOLHPlnBBj51CxwsvDUtaogiot/9Z4YVOtpZ+MEhv6K
Yt7XTEUJf8fdZzqDZUs3lmFFyEl+80YxpqWBBDoMlTw9JN1ri0ZkrAi3pUkxbw7UVJ/NcAgJtPwZ
oJYKgmgMrClIK+1G8UAtTT+7k/+8Y4l2xZZ/J3Viywd/QloduEWU/VoBfzdZZaycDS9XB+quZDz4
cYVI0FfYpWtl5FY4D5odipaI6jSGxsUus1I8TR1QoppynTsO7NHvVw1HbqQhbr9LKed7oNrWCF7z
P6G+5Sg0sCHJY7hnveSUjFBneRKMlSwVG2/Vrz+qLLqGKYI2/ce4ObkJEPj5eHqi4UgDzDEYDYVm
6gQzReYfFiV16J3F4hZcVTxwPQ4WAhZEzpDbyepqbUcjjnQdmvxjE3kYaPtw8wZ5MPjio0kRPuJV
ORfZ7LDK0F/zbf3Y7J3cIystCeVTtS+LzI4Gxw/vv49HLNEgQmV+L1a75XStfB3ZkFhDKglOVWax
wYEIKRcs7khQxEUTxc5RJ9htH3WLiyC1O+U5dJuWjkC0Kx8HBhA6cyoueoF/GvqjRlZB2xlAq0ED
bula7UQxtd3/9yWCSlzloPs4YZZFuNQCKvHGT2XVjGKaBXaYB4VfHHM8fzR9kGag8dFcZ9Gb37Nu
EGYqKVZBfBcQA3HbbbAhKa1q8iSvpchhXmokduOW+0TvY/mEgSQaBZLn3e6qYfVh0PBtRCemYyOr
b2AWEIpzriOdrlF0SQQPyPopU1hvuUKKUt5ayGInbE2MIxbzEtiEJjdrZZgxdNMDDAuu7QQRL2ac
D0r0JcIhFwkOQCAhtDTwW4auEoiJEPyajWz/xuZEJZuBZJ07PnShTmoiJGvdvpbxYcfIwN0EzSse
hd8zO9LWY2d8uMXAjUgBUMudNWmlbv1sNnOi8tbWCH0E8OX8AgnmIKmyMkU7swZ1xUxIwdj1II2N
elrboMS6X4Sa+AP0ClVv2ShSi7ZMAFapIuJKvfOm6Sn9QZb8DXLUbs+J4Qd0OYuCLC+SXDSLUXi5
aVnL8wyEdB/XvLECfgxyUyzwCZSippxiCWEVqPZ3vA3ofN7NmWnFNTAAYYadd7NFTid8x3TvH0Nt
ZqK9z6vdNWGEuoGasgVnccIsjrRR3Bnw5qlWv+hCNvm+tT5uTPK+Ih9ualI0AE80KY5aKWNucErP
BbCXb6FxjtWO7jq20z4QT1+wGNe3019r40G3zcnTl+k4EjoArukUps4tYez1ic2hUx/B9y2iuKfV
xBRuv9toztBd4j0kc5DP6ezzOLgwiwErNW3xhj2Gcz0ViDVrANoCvwJuIGYSdDJep+gO/wWev9f5
rBrhp7PQQ3wlmFh8sFhbL0E6tpNn+KRZp2PwhDLvHQLbt4/fhLe0K1+BHIoJvphqnwTzTHE5hfw9
ZLrPGx7eWhXTlFC/n3e48ev7PINIAyVN5icn16sZROtV95Y1loflf+czJZaPN0rE1ZkhuZDVWM+E
o3S4BPcd5t7YMPCF/iZG9b8dPlOKKu4q52hjZN89KxFinTC7auP5cyArG6UnfHcKHBkFOqoVvy9L
Gh3u03OlbmZl/ptbozppiiEv29Mcs31oR6xQoieOzw3zPYii5jkrVNIe5mUEJTXTMwbbECx41TgU
74aeed6CDIWqHXgSO1juXFeudodFDLKEAvnJVQ4GPe5Qcs/zMn2s1q4kFW7sLEhY6ujjyAdayIQf
6AxIsGdhkr6iTvIamB6gu6NrPerhGAnc/9EK+I3NMfBh2n05pU+/5fPiSlaZkM2bzGG+tpJ5rHca
fwko//8CXnycn8v4uMxV/iWfy5mvxDtjaniyB0jnhYHq762sBYQsShHc15WrY0nBGBKMf4lMwprL
d2Xqw81ZP6Su8K8h+E/fSmd1sg3X4OyWcadMK3KNdpwWwBlkvdqPaaZLE5g6Gj3HI+3nFfBPzhNA
3NJUSUZn7cYnZ2n98SHxZ+8nfPeAdwUYREWxLbrpJqIXSO46BiwY1gpoX7yjJ/gdJ3rKqFCsSsYo
CkewgfQbBtXKm41nJn3WpOKYec1ffNM+SamiEvAhuE88Dvlmtcwa4iJmTOZma2hnG5L1A6qZuUN/
CwLdmaMVbOyu24/5SHlT8g1StZ8DBUP/Zl7JQ0CjhsyufEzyHgWtlikWMefO0TrHqAeGWJ1006HL
gstTlNMtoNKtUlDAD9mmgynwHYo4EcCuxFgQ67su8MKMJ/hhDsQABBORC8suVMqbo8Zk6utvh82e
wnu6mRXhll0cbsqdZgIHBHes/b+wcjP9MU10A7t+Z86VgBzYP1D4x0ew+4yQgtIja//BMbV1sqLK
kBktboLdgFKIAinl70bABHuZytDeZyOz+qv4oJLHlRiLAAHEYjppiT/lnbjM6z4E6RDHyptxN6ju
Sj7cm4MdJiz56zi9MM2NTR8WUwT0nshJlB+Wp2Noru+4Icuf6OE9fFeEz2ZLMXNclf5bR9WpfnMi
qoCrMUPVX5e42yxZ3rNtdyTqbBk9om7PmcKJQDEmKM7MXWed3aVovDSG2RmIrJpvlDFO5fisYuwh
kxZMuH4RaX5dY2XaZj76leoEsumSOarjFAnUgDPjuhempdyD9GEgeSIq3RQM4PYdPaLzhx6YdUOo
+CLU191KW9c4Rmu6R8xJNVQdl+/wqwtHLHlut6gpBvFXJw1F0HVRzh6zIgr3nu7pLNkHYC8RPtjv
Gtzw6+cY1yzPQXHbgBRR49bfcF3dUdwggwMjSPBk2R/awODDlQIILbEOAG/tzSkDpivdS9xPNeMD
tzGR0pcd3fW3wXs8z6VgKBRjDkjWmNn3J8sG+MSBXBzQPxi9loq9K15DWCA8tcCditGEFIVyeJ4i
mghTljM/GmX+DDusZXHlOzHVcHNBWBAXAhI0kX3/f7Sw7RSFGHAPRMi2qk7Xaw75AwjQX+XRws+j
B9siCQGHy6oZUjHx6KK+cp4Cm9tKN26V+a6ar3jSbRO5ig5J5nFfjD0VipUImLbwjkdNVt8x79Es
/8b/5vLBcPCwy6ZcWxHAYdGzPOONVlUZ0uLG6GaJFXrAsAkgqQSElLmI/BR/EKD1ncmcmGSWdIBq
9dicCP5nPBnPm1rOxLKT5a903YUObaAQ+cW2hcOWA2Dgr4PGyAlNL2ECEEq2oLp845ILncQRJIW4
iAwfMjwQTK2j14AXwpWMqYoFaFpAAD8me1hsNuMV5hW2WHpzSNtFQn/cWHLsEkQ3zUhyriXfhEdZ
RM0rsF8suOVDNduX9Y4KT3E+UyGkBnGwmFAz2JF1oUDISfHKQlwzgeENt7hKcaQ5MrvWC+KaQHGW
npGvHeVqPDLLWnf4nUJtq26kJx3t0cFvVzk0QaNhvZOjdyXscMy6u2RW6K3jezLjNYMK/AwpADKH
5bn/i3irQZKpfVkT03Re8EhVpgbLoHLjK441lmGEx9WbIW+O5JsXEeqiEYE4SjKb9sRwhgepiAVx
moYbwIslv2RK4kMHMNrOh9rIxMRjxRGBOeJSTPZfjpkR8F2A+XZeTQlnc2orBpFc38qQuV/Eyyem
V83mhClXxabfautr12mslC19M06/DMMNeCGliP3EP6c+DuIeHYGGKhxTaZ6QVsC5Aj0lg7SduHBf
ONrcI+qdb1HSzmLXh4zF+mgrHCCfkeYjLZ1TClaZ41Wlry33DMRImlO0diANf2+oPAkwBynZgpNa
06V2m7dhh9StG3gWZ933kaigAwD+E86Vqna+GEpb0c1mgkyrSSV9qXRWowPNv5Tp3lVNTwpVXqXp
WQpygSeOPzuxLS5mVVs80lpMjxM95V3KLp9DHbARa9wWgEdD420tMYVXK9SgEYnH/VHHn+rUUxpC
FYw0zV1BoSmwDtHfxixvnB5yKJIxD3wIJrXn5Dz8uSy/+C4fI2/9SprK1AKJI4LDP6NdYfRwBsGj
jzmzGC/svA8zzB7h0b/dIg+ERQOOAi+8gBPs5JidbY+x8qk9Cja7sHD7vPxJmuaeXEqhy7FSu3Rm
f+US2YzTV60vUlZ2ykPC5UfZIrhGNh3PTWCNFOcK8xSrcWS8dExtQuAIol+J4acU9FyEOU8PYm8b
LLLwOmHEo7ZFjbTHux++wSwl0Wqt7ivCQKwC+Ms6NBKawMZL5SXuLp85rZkhs09RWRQtOii78I56
u6pst2aXCW4Mu76ZL6EJH/i5FIMe0RZtvvueXPHaOvj04of2c38I3PH6/FY1gl1Vh+iKhAo1T7Gd
7q1NPGKeDN1WcxumQTCcuaweoxtX0/SnFFVwlNAbrfPVynXlE6R0EwenzpO/PJCXvPY/xScB2S56
uycUPpY/NuHrvlskDYEH/TuctZwoGkp3Ar539qLURg7E73jbf0tatVIwZTUrSPIgvTxsy5JGhm3f
TzIk+UlyC6LVm6CJhhlg14gro7OfQVvRu2KmH2RTelltSm2zZmskGNq5V6mS1SdVST8JXFTmuTQJ
DOG+jHjTLiXb1ji468LvYiSHC1cxIOr3Rs18epoRye8hFL/h7xZCP9sbp27Lbp9x5hxRW/4d6KX9
TK86CqgH6S6HKBlaiGxX6bOz2jApimYrEv9zYWtYaFVUCDBL6yZ5yLiDavQuTjD7aVz0lbW+/LHH
FBE2HbFg5yT678VRpfxQ7Klgiii4UZJ/XMBBQQi/PnrZmifTTOAvxOOKB49nhssruZvPBgg44Ifu
XH+RSwByilyDBgTOLeofekqWaPa4ASvp0lsuVx0jCVbsmnIY7aNk0lpR7QFV5WMiSdm7cHK8YFwz
vszxvo80MPBi1i+rBvMAdjcvweQRD260JzcQIj9SYuW+IHPf/eaYQb6hOmAdYQ2ugrZssUybH1SF
e1PAw/vDU8LMnPVd9UjvfSCFwXCt7XFw57jVsk3B/iLZjrpjQ2W26AxMxYWP2MJkro6F1Ea8lYmz
uiNQixYQ3XztWogux1fyCAjQd7d8BXbzk97/YRpMMwtAcwHVtELaKENLDT1SigxmpF9DtxF3cC3B
Qwp0bvTotlsBqHsJg5smgZWOvuSt1ss3K2cAhcDHtlq08yZRSKRNLV+vSSn4FaVCq6ezen9WCO3S
B/PHIJ/kKMIc+l7CC7k6YEKu+sczFwbRGOlg+2RC9zmx2+t5tDI3U/ojahMYtIt4OWN/saEFDY9M
/48jET4vsdUAWX8f1jva2hLRs46v9Hrwdi7+0QZN8cAVcU+yn6PPSpgvWBG7olDr/MjKd5BNiKW0
Q3MzLNVkHdmP0/bmWL73i3TgBoylMP5PuADZOql76x4PkpVNLzuueHB73FXBi3OUw9Ms9K3cxxsw
f7me6dtmL7Qx9lsCFn0l6m5jO4pp5xrbcEUBIU0QarO0OOkC/Ty58M1A5P0AnyL9SFyoj9/gTYKP
xd184H3PSzypuARM3fJGyBIH4YG+eoUZMpxWHn1FjQ5vRsSPIwcFcBuG77X7c3fH7gen2y9Q2id8
UoAe3S4m2+8TdTBuwcDJxBKXcB5i7MNKXa4LmnmN5ghWg4MGyukMwspf5vYsqhyknfGj1rRUNoqM
HC3RJAanNEpRG7a70fUrbnP662PMcpE2GBS5RGCMqJFwwRbVZ+moClFl2rusXTUTWXAzVkpGjlB+
e2YcTY4l2cO/bMdkQ6fBpeSnkxpTZyd7AgPoJOSHetQ167g4zYQeIVm5C6PirS/mn+z+Jl3J7gVE
Jj7s3JVWgJdjuwUSc5qvVrvDqdsbPp2Gy7XIxF+LmzHcgdTUyIaoFWki2ufZ75jl458cH/yOXJqc
/EVs8GIhQiJ6vZCprP++GRBYPqomzgayVbLgl+NTvS8HqlZ8ItCg/sG1o/hUcIx7hn2ASBA4MU1g
ecS/YfnmCUz+2MIgIAhyHjRuWExTF+2fegq6sb+SJQZlXv6glARH7GWLBQGL/o0bsg6Kn3aQcXO1
4MAKo/lCBavBaBX6PR6FFOlRVwqNrm2Rtr2f61YYrz1c2/YXE0IbOPnE1wLtCbq4KDj9vvj5oA2X
LQQi87T7yxil6yLKqEhbcxR1NK0k7QMs2ZqsUYt42eXE8N6e9eMaRkl9nQolaqDFSdmfz4B+8fDu
ZMFZ/UR/sz16YkxZIm4dgjTT7ZQ6AG+/g4JHKgr+LGNUnqmAJHUCIHP1nQ3iug443DEiM5eL2FmX
409KeXO/AFJsP+NxKByLga3T0HcnxFWY6vq7OwR/WRu3+gPBkfxdMW6nNuqcuQVibYm+/j8Rcis+
l35XnoMTdjVFDNXc2Ji220Hd2ZJD1rSv8i/ZlMV1sgnm2QhbRUJyEYg2VY8bFlezxg2dbFwuYy7A
G2U72u3n1WIrIsto4jL3fxnAfaFssivTjwG+NF7Oh3vrw/8aYIblbdfLociE1KJ5+jmDii1nJ2Kn
rmGWfJd/0PVF7Z+WQCiPEfAsuWaJhbx2azDAhmu+CDZNG5BNQ882r8g4MZGRvhhJIpBwyOVKKa73
3wm1etalHZQJAr665wvUjMqdrFXqMH5hus8oBOUPzqypSdimkwdeS+lFekV+upJmJYj22RvvszTY
4G2nbK8/M14/ilsZMMCOI6cr6NIB9E2iEc3tv1+eC461pgrSjwZ//iEdZLnGdcAAUX1EbfOZGH7j
JKeTsxti+PthS5Aj0+uR86gt6z+isMBV04D7A+8Kp/IihWZnl9MLL55Rfn/+Bzuh9H44xqLMgGcu
s38Jt90cG6Dm6lvFN2aeSXPiqqEhgv29CeSBt0RmVX4bKYxx7/DPvADmBDwzssMuEr4m5xuEDobs
b+4XER8SsFuqroulmTZJiUw9UQq2t79Ih9xq0oRsTlxN0ku8ImX9D5w3Iu+yrN927mSzV9qcjn5h
NFd60IAkZtD28VAiaDC/ciAI4XQJ/qvwC9DDJT7j6Ek2ljil+EnPd4iq5QOecMAAdtktgdjIs1Oq
GW0CrYNPhfvSKIRTkmopXKM5xDlniHrBWZG6VIr15z+w5Z5IRcRxrgj85Wt3xjLb4+TAWUs5A+LM
5bm/8nn8VfUFZjvo3Ak2qevx6c+761C96/3pNlu937D7SGTeCHUeS5qFzjTbP//6iLVkoZj+/Sue
VoEDashSx5XZ+SuDDyvFLb5ginDbcxEPLlHGhw39VtkDFPjS2nsBHsnjdD8Vkxqp4EkgHjpnoly9
IHCwjKCBtxdII883Xch36LssuHpDyU1HloQOSY3uFUYgEs3Ym9OPKxET+n+xbICrTg2OKNHHCOEJ
xPK89YvK1nRG0tdxde0S0WiwV01jJJ1RqegIe9GGFbecG7UFruH/yRUenLM8ncniuUhphBrrgy20
YDwfnyxwQfagkmUQbK2sYf/jBxV7i99lgKnbZfkwARiuG51ETDVAB05dKFbke16uu5oSFX9+Sr1G
1OVs7m+sAjTihoPKK4Jhzb2rKEyFkVtu66ZOL3hL0PSBOiMC24BsNKguCtzzV0QpxjzOs+8AVbYH
IHSLiLfWDzMov5TW6DEg2HshvO6iTETRGh46kBZOho5p4aK0TG7/9Deoh5ZKU6T90Qm+uh0Lpt/9
lhF5QGrYdjIwzlNDiljXe5Jj9lOd0gOMXzFDdex0Us8XIIGVhTugCZPm/2ePEdAdxx8/6rQdtIO7
PQEFXsj4/fY1Ent0xzd6qeOAxrGArarmnV0NMI2msgs6UdKfdLww68+dm7H0puiNaoNpC3ffQ/YI
+TzByfRqaCnD5ZsfqTahYb0s/l8M2OAUDioXtnHmNCo8ZB/OTxpH2s45N/Mp6qkQt1GKCZVZfbWC
f9SgxIAmJZoa0e5y0dJz0GpCwS0qBnN+OcpXdDTCoEpOw1ezX+ObK8TcyiGx2yvy7mO+cF+ofkGf
giFpjKvAbTqZZT29/CF6uhIa1Hba/2qkpubwvxYSPROAwHehA12w6iIaKH6f6sbxlUSEgHJQaY/O
UK3n/g/UYdNCjqpkf49mmIz/AQa9v6xYTmWHmHuOlzDQuvn/rC2FWbAluvWV6qjofQknKA3gEJjA
y+MoUhokxFL2h5K00bFO845WZ03TyItlXa/MWKkInikELTr3DcO85Xec50nSveiplHVVu7LaacQx
T0QTYLvpGV29LwUbNR5UZU0gFkzoGlz0dm2RIH5Q0FJhhyjOJBwc98gHYqMoJK2n7xOiE5/670ZA
/2ljVMli7l8qlvnQYHr5uD3OpfWxi8t8iYY40R6wQ9RS6UeBhRxV3VC/x0gXKTq+TV0O+ydmsgKG
/4OQ39Vaq75k9jrbCN+jc5tD/SayCJfsrNeY0SacYes4xc+wCB9SwwvAEZtbKAUMYqkCk9Y28CeD
fIVRmASFkxI7i69xAMm8vq5p2wRY/GkEoNV3IF5xbMX8MB2jdsmaLeS3jcAk8ZxHEKTT+vRUmbNm
yS6jNA4YUiTg3dOglQDNqNJXIepJ2yRAeQFn0IZxXSucYgVxsZpN2Ogbr/helqMo3MnFA2jQu0Wq
C1SwoXDZh9W8dlW6je2iXhPw4EFbOKIYfyhL3KVqtjUMVG5i3Hs6JrcTRKADKrsuqahd6lsk21vB
0BIWgZOLeV+RcKldvVpTl5aYcrDuEaAaNFc5snt2dXYEsqVgi2yqJ7IBhdR75vSBSLvnlHFwlV4X
zkxtU0By0eiM0NK1a5gV/ygnVnz+ySuBJjw5crCHN8RBKH908GNCt8ur97u+cbQxn2sFCsFUQ1ga
bwWIprabJ8nfN1WUrHadosLFOPgMIEGuqf6uKOOl1RhA7K9QKkkiDxir+lWhgc7UqYJl3HmATKJP
aGY6mWXXWmcz3e76PqZzyDd8GN/snODVzJsKyQRwf25kNwP53kRp64mrhCeodnqDSht791U0VCHM
2xZgrgX/BvvM86ZRcV+5WmeqLyQzqFVLuYKWO9nYrM+Jt/sFly1tY0fqKtzUkcc6OmTfm2RRa7cP
ZkCzBbMkI2aOhkyxyHtWgH7HSEDgzCs4afRAWCae3JmNzZavYTNy77MVf1tX86+68oxlnipj7cod
lM76iFloZJ2HPoaZMqgYT2vdpnfRMD2bXV9f/CXlkBBCZxWHcRbtpbRx6ynYw0ibZIyK/VsgRF1Z
FUZA639DukArzSuMD668xFHfD5OXBwQvIc56cvIS9lgf3egIlqTJ4iDM6iJW7rcvE+N+IfVJzIm1
nwDfoqZ9cuDXbSLBt7ZiBSSkkihESGHfPSrGqh0TFWRbY7wiQEboirW2y+EdOihxLn22sneu+2RL
SK0Q5daJFI97mAY4doSGmTs+r6RwkKvnvHyj5jxqaEzC+0j8Mxyc75+i+lQ+G0a1OLnbdl5Yy7jf
FzqhCGLFVM8e8ADcn8jTbQGS0asxtTh2NeDLi2oY1THJR0Y69Ye/MhZLIXI+8vMJ5fVnC27/i9Iy
Z6GrUtTpMsQPwhqMRXOyl+L8nZKB6M2g3+O+gDkVAQpQcP0PnLimSVR23pMjHDZ5V/m+ju4Dni0x
K6l7sSqLmbGw57aeJZvWeuo3A8vvyg3RZ9bmBH4sPZuMzjUoBv9Kae3qEQZvgNfUynkk0Kg6U/J3
e1ZIWuUXqEGB7e+NgVH9cmGytUAQbZLKUEST1Yi2A/TfR2+VQoHdJyny+9xHJ7WgTM56ODk3nwua
+gnDxvm1vio+hFQt8C+eq7E4qcQV8QkuNJ70V/Xg9nY2tTOKLxYYfHFgzK4gn63vdLRjdUJ+mHfN
Grpv2xm5HfdvAzGZCfv8bUtbKg+IW57SJQl+DD4PAowveYc1bMrjfLs0Nqu2mldSAwZEiJQJzVjC
r28E4job2vLRgw+vNIJgL6yn/g14q7uFniz5cGwYbEvLJVFparx7dfyBW8aWt+naQycc5GQWrcE/
u42Qv5DiV2js53Lf0bteRDldwE0P7RwEuTjqNEyEfOHk73sGXRXByO7sxZu2Uxw+VIb62xoUVxJ1
msrpnwn0RsiRllm5IMpWbEXjv/mG7THcDudcGok9l6LtyEQFG/7Qs89hEWX6R/oBAKU8yvZYG8Hq
r1o4nQCX8W0CNPqcI5oNjMQx7xbl5IB2bsB00Q5tAJRgB0b7U7wFxQwnW/fHYmH+66vkh2IV3jzd
XqUGChS/zAg2M3OuCXtgycArEMIl8M6ncyvg2D3DQmFkKcNdU7P7QicGRi4cwu3eD3x7Mw65gXOc
+mOogp8ksBsf4VgiEbsstoiM2wkHoLsgtbawwL4wJCD1tlx6WfFZoFewXAef5mUVsjBocfBTiO6T
MmStXAVc1yrnAfDUXooDUIpayreF3oaSSDHcpiqsVRyDzDa+2T5tJZyfwgGfHd+J2uYROLr+OcBX
2LfPVNDgc7OFKVc1x+srOJa/0DFLBwqqd7+aYLs/cVuCTLu5kTE/MtM/48sr7RUJLLcfhIo2IQII
MRrV5sXsVugH1j6/PXDmVH2MBTEwvVEB+KnNRRwMW59aYRyG8kDglCyExbszlw1E1S4GJt1SR5dQ
kmdi115xTXT9evnocWvkfiEP7XAcVG6qXN7NUqEqBimkGxCvG3hydH17nARhD18C9wthvHjQK/wN
Kg5gpY4TSfp0bbVnny2574B4lr/S8+D/WdfBHmucf6IlUzdtZRX8Zn+T4y2IHb9mk1nwUqBlqsfi
u1cO2JN8b5lDANLAZUMIotp8W0qEyhX6mlNAVZJuETtcBwq/0eyNUFK16FR6LjT023GQWixXDH6f
6mwnVY15dRZdMblYCo/fiVz5rqfSollBdcxWGMix1ARwLhIbSVobGnF+wBDlMhITowi7BQTp9ZHY
aO0B5CEJVIqIIqadp71+gU2hMV/p09Sl9G1wX1aMUmOsX4aBp24gBeeK3dYvG36gpZL8TAhETXZV
z9hsflSbFQ7hkCDj6o3Yg/6542nAv6beA0kDbOrYzVRUFP41xEGGGs7ZRpDtwzVSr7nzrXEV8Jwp
7QgI5FWKIOEpJfHKbto/hXANWt30ehqNgqGppCPn3c2R/ZVx86ThXv7Rv2SLaY5fdzu6oilHa9Eh
k0ufG+NujN8pOrzbiK+/Npu8eL3Z5Mr1B+tKygyxYDhfx/XKAWcd55EhC07IIq6VNsLiQ0CLZ91u
b5TUuHSgP3X8kQthh1hQJBqWU/9wdvjB97mu8dN8rFjChIGFvdVswddHZJJgRmCn7BA8wytdKD+n
C23ZuFPq9XMbXy4rNrKnTIE/6ytAz4x6QuiSIk6Zg3BKkUdFi6amPwgeQh3XpkFK7wDFrg3a6GTQ
qD0gBLvG99Db36c827ESEgId+yS+EeNCKACwLILqbOeesMEbN9HiMh1wDO/dTGquGAe2ljT9HxNn
nIgxY6KI9XD9eNfy6oE/TQuJP+JygLb1NRxdMgkhBWCs0xC8FKVSsgxjd9g77b20s93Dsb0smYgC
inroWJvRqWPBVZUQvLRNsKC7Vrs4Zw1MCGAdMaXTYolUD6TrU3t8OCN2BievH2WzPs7i0cS/dZql
xr/VWCpXdzkiIlZwzXeZxnqFyAyfvQSym9e46Tc/y+7QSySpH2k/cJ42Ip4MC0G2tgpHGejUTfCl
0iGwNYgzeC09xBuVUHJo9xbqDDA7J4PmfuCjUU2uBVv3NMnd7WVXFWi3sBhF5q8DnDexj46CAn2i
kMqXTHBncDI1r+Q9qBUwZWPUcDbLcMC0o69E+GwSrLQ5HXzxo4ruEwuybizuXd/m9SYNM3K/tyuy
t98AXTJdJM2euub+XJ68fI1OUyT4M2cU+d+hmDDouZGGaLPx2r4GG7yI1hqAA+o+24Dgq9O2YcU3
ynwH9DPIBwS1a7DEGp1C4NXMT8Dl68hHYID5dBgqL2qgw+LTcF985AVSw45926vflFKapmTVdhvm
PoBC488WSDTDYIkxFjWpiD3VaQmCbrEq/36P/anZ0LWOwYhctSPSFPAKcAnhZDLk+cMNY4UP6mMM
GfWAclADC5Fj7OkqiqNiTLYHx0GhmGIrmxhGjGburpc3qwuMfu4wee65LiXvLNtV8wjWF22H6EX7
EWkAXiNx/w0E+1hlQqQ+I+J9+xV7qQ5nyWutm1VyCbIXVzKdHAUDAGtqoHe71wrBpWd54HAwIYCL
DJQvUf6iuh+6Ff2tA4w7K1pJA4A2MuFAJ7/y4juFgCp921Gbvo7W0D8GKpXFkci0WkC22jrPqWO3
Wi9XHor7Rb9pAW9ovmjkn8lqlYFNd/ZYu6l3kAI5oPO3w7mYHlv6vmmtAIZBaf6QRLbDkNJU/XHv
rc7i0TGdY+fhSLUC08JcvNIGw2bBxizcVvKAEzt+zzVlc9NCAYQL8nyUlI8UWIai1+12h6lTJ1GI
YuJIxwoI0x18c285Z3yk2FCqVv0cY4tXMJf14xKgIZMyZPnssdu21yMs7qsd7fpKqWLeJ0FG49Iq
K1pdZkPA422UtaWePywa5N8fsm+XzKIzj9VuI1d3OlGYha/fFPCch61KOi9LuU+mxI/w1ld2pXQ+
a2FZaOg1UQLcdmAbdQQlub7cEJoaJt66SpuAfEal/zvQiS+iQ+mcWMBtVEkiG37QVXMF1RrWV/c6
F+jLn5o3SB1UN0xdoFH3cXJ1+PesculDJmaX2SO99P6jFkpqJfmGWeYL9I1GckmP6KeZigL+TEUb
WEZYfDCmkB/lcc3LZccuRFrzbzwm0Vjvw48PMxeprIA2tdrUV3cuep7hgE0aI4HbtEeC4Kmq+YG4
jjzUSds7jQtXhaJ1d9GIql7cl+dAktIITy3ZzWpJIIYIO7N9LD1WAiDPzYOnFT1Bdniwn/32Y+NV
jIEQ5qLFmAGhEfdv2Wn0waLhGc19VWtUsu1CH1BbfdIkAwJD0laQGvW00iLDMZ0lBMHSMyJ9kN0C
KwDP6h17fWPkz/sALFbPJe86xbUxiGADIzZjw3TWeNgMVRedHATss9oC5YXnxV5uVyBtJwjSoX7T
YaRGu1twUS/MJbr8t2z7hjSAk45C9eujeMlSO95kAHRAfWL7L3rR3njus2Rixi+Zxv26LS4zaSua
b+8VvIzZ59/tpXmCTasAFw4/+0bYNT/JpzHVKdlanXbm+EW29W6End9JfMxaVCDtGaZxx+9SXALP
gU/VyRLo1zQUqD/Y6o1DKfIY6y/EagNWhhFPXTKS2sk5Zf3sYJ06WFwPZfoFC73xzuRvs11v6GNm
w+wJNEg2E5r/XtbRYj+TMRzM6MtGcapKywPrbXeU+UEX2MjqKL45SwdxV9WdlsfyypJFEEtZnXgU
H7Aho2z3i1JqAPUUKAq7XGyE2fmzyOCOCbC2lxVsTsyNGZLH8U5jOyXdtK+j9rIKaAReTP8mpyq3
6DOP97T9E3P326WGA8mV8qSTnBlc0wixzNc0BI+Rvp52tIjsUDE10tTK2kSOkpYPbrcFNav3kzGP
wSWEN4wUCaXzAyiMpihDoeAceoYdI7idEnfO4xWsLC+aF4lKoqqxZR373iFyuouhCJMv4Yf0naMr
+GD9zrSxmehsfUAdKo4OYKUDnnp+imH9/qAlBy7jTKYK37GjOo8OkQhLRtzShQj0PgZBdYvhQjKK
sqj/7wD9o4niIdnCiQhto9uq6Q3gbz2I2+9tuYvvo2d5v3Nw8/UhaWSQYLQDxy537BKCvCAuIOVP
Wtv9uiythbjljvDQQP33sdsueORfSpwSwN8J34XDcxNXHp186z0Zk9JU5MT0ia82Am710ZjUbW8n
w8sj3JKZhe/pNkPXlrOFmS7JymmGhNcvB+/XwaPUTMlXUhM0gIMRxBDp9lP8R+6DPaQOdUBnX8BC
X5cjc6xay2zhw4TTmM0kdu1T+ER+0PGvrJeUC2aK0RKc6KumMlXnm45VVFH0cUOMRUtHNp+A/F9m
ZJhG7siTnH4h2BZQtnQ/LL7xReJQ4NL77OWsS3/ln1mxCYd8gxzKe9mrTPMbIN3tV5ZCVoimQREd
Ur+rY5WoJwMhqshndVufvCE7M+H2+S/k+BhRAXfr4RwBPMGKFitdurmdHlOY+io/jPy4ui3pleGq
zpDlgpln4zKBQqb5heqtgP2GYQUq7Mb+mLb1g06aqUuCO060ivetHjlpBK22Lo3Et0SBUdXyiBc1
ckTGLfZHpcEJcYQSheGyoVWJ/WqAXarn204vb9CFkOT2ToHeTdWOgWUryhsUv8HEbbMv5hUybc9A
oaimMbR3EbogO/pYvILgkmRQBcLXzqGcuolCNPvc7gw5IMFDbgTe4qNo5vPOkQVWjn7FxUunZMJL
Z6UoOcKLOQsoiVENi9xhYUIDO8R9e0ivI6MkZZHIHzygfz/QyhiONrxayX9UtxHwvnoWS48Wvl5p
nmipLUFFzab58okNwqlMbuDCWVLPuIuJY+h2lVQJJ38ZY+PRmICOn1FJcoqf1b6FxueCfi1zNkli
shXhLadD1n8+Tbm3WHP4gIp3FJcT0RBvpGUDYV8HW4Q1Uzja/ftgJBFjVVhhd+L4PQmeOe7utmnJ
c7emSZqyuKcpW26/CuCBPbqBIEHRg6CfphPcRJrHSKJOv/0Ar8x9B1oe0CHcLmLVRIEQl1yxLiFs
bq67FRVksMsbtVfpYyMlyksh+/tDe8thBH0hGF5v9+4cDJ6EzMwE/LijxXVIkwxbLX23/Ot0OYk3
xMqQWxmzy8C7nxOOcjN+21f8kxFp/93KT+ZuMtHdUcCmRyerAJ1i2HwlWBQMhDfJqcaHgpFP31yS
TwQmR+nP+yh4UZ1IovPGiT+0J58T4LQbXnubbXW96sFeHaP/FORlpHBSseelVsWxRk2NNUqqM+TI
R4PsedXslMHMg3iHvYJSdwTwflEoNC4GGGbs5DzCxeADd8AhBqFpqUI+kivo2mSCXRMfd/oBxU9E
uZ9sXSr2UVZ88TP3mD7o4WFhevTfBIhgH0GwLUFDHtdPYgN2YP4r7WsLYN5XTnFDMvAypANEm+0Y
s+8Uc+woCiSrYiOFJiQx3uFylVmeNQae2f348DSV7QrBenHaBKzc+vWLwN3AysHHFb2t1ek5NBTP
4HdRahBg8qRYFYUxVGwc/GajGkWVn4IQE7kgPmqSJd0t08yN2mzk54zmabg4EzlFi4tbT0416b2x
H2dcGSUnQ+UCkiuqP43/57W40fyw45CI563a2H/nveYOuGYLFKm8SzVmlfOvN9GtPnRxXbZ23dZG
geQ58sONkgZwf/PvjRbSxnzteMMCriNK+3hxzI0ytiABpl6VVfVQzgR5foobLg4AfvrqqXpe9p/D
MxynFFJmzPXLMl9CBcGbcVoz/stYas1u9mM5xEz2ydQuajRrCAGlvx+Zxj6HiIAOeqQo3FZhsRIR
rzbNfxksgHgjsAlmLOjmJGdzX3cLsyUpad/bp19kOJ98S1D/bUdHD5Svl0jWeSWrQW2rVGOk3NSq
CXeqio4K79X0AIIzAiSm4J7o9wHFMO14pUT+Lj8Upk55RwHmGPr/3mlne76VRQMRXPt0jFg/XAE5
xikkQBB56GU82xjLQA0JLU5ZhN4FnLb7NcRXbvNczuZnVHCUn1h/qMp6ZaK1J7IuoKRTHeC2tIKq
+u2ECe7ucw0XKvX/mCOJefxNdz/F26xfpjY+jPTsmE+tWNSalO7acIln/IQin2WgJ/ps35aWh+n7
z2809ugaztpFUEGB+VyEZos5dd3dqlYL2MHCwRHwh3XQSx2AqPRPX5tP+u+e5XnfOV7D22661Aos
oe4jFnWTChPo7KDlqMIry08EbyoEJl+gwNOEEz4LI9HQxtoraMw+wl8rjBdyZ1vRyLXGk8iT52pA
eGhGGCBMA2oPt529TlGzvpDS8cqVmOhrbUZbyNvY4UbYX1+Q5wwHf4qSifv6t1mtpsGknmECcbVF
zdhfy3Xququ97pc6JG/4JBNtnEhsMCo9S5dCfu4KWpeanIhmlGIwUDLfR4cAbPr04q+VMOIx5T4G
lM5rvZ64E9xqUXH7NEjWaBCUS0yIuLPuetd94BYbRE4F1wldyaaZmWVH5JlziGWTf94OW+XjL9E5
U5kxXL5/ueDt4P1/FaAdhi/E3gX+ykQVi79WzAKTXhXpN4JreSWtXNhpRqDI75ei6N7XCi2YZdc4
z1+jtvtPhY7ZPvfzILyUr6sidvtt/DO8r4+HdP3B/NNffnZdA+6gQxBZyWCJS/myLIujvU+Or5hQ
JuZIHe4ycLs3Esx9kkM/uVOq+YoNM65APfnfbwNiQKDdFs8zKhNWXBn1wqjwqz+DyNtA1SwNGU7c
/y1Mu/YGuoLtduA1XHLIo9w9BDDR6/iSyJ6mWEv/wQb/1QoIEUA+oA8AvJXhYFy0P3DKYM90Ak74
Z36OGp0czjeUAeiE9/If9RVLxHw3MbtGmwWLAgK1SwZivOLeuvfOnTClB2KSe+mS0/ap04a6iNwN
wVJ0rh/o7Xkay3gy0BLWofZYy1RBy7OIxVBzM0P3gqnJIIEm0Slr6suTtrCoz0im+Ko0VLqR+uxX
vIl1WEa70XF9owlUTpVa8XadOdruPguLQViRxlOtFf4rjU9PxBIS65Hy6hv/8bPTZsxVjlpMgwWm
CNH+GkTPPxr9koTcn7o9NWqWSBQ5nbKHc81NXTU2pATnr2tAwyfGxQ+IxofxVXIemXNUJK2Jyxhw
wpCEcmfZrZSZ1/ELAqiv5FY0cgJZ//IPvHZMCT3tptAoEDMbcJfaIpQBCFYHKGervWtSMThH0oVI
z94hfp41JZjcsI+tjMB5bkvdgRjY40W7UJWjpHPqhCgMkAK9xYClWrCMcSNLAz5LxjMQKoT+ywE/
ulNemvFS+5t2RcR6UYCO4MUbRBkEMHgg8M5m81azN7hiSLglzAB144US0gkSMLQthNps/y5i+oCL
BXWWFYeYlHcGe8YmD6cH6dnwCitfhVw7FalImFwKun5u2TGJ4bJBgCtp568AGPpPeaAkOoH9PBEd
0wjROB+X+1ayttQB3jmN/o1K0dtDDfn/6MgfXMisOsTNV6seb7VaJu9QUH5g7E16zJyyHoZ40M7r
U4VahxXdltGeoprQOIVrUbF3eQqJHk3ZYB1whBpPyc4S6HPDGlToOt6IBmEQVujXcibOyaEt64nS
eTLRbwvwHl/rsvvWJ2Y+7THUhkyNX4+RTy6UEcReIHFkCOyb7MXLXJWQl2XWi+4zmZg37cfHlm86
6nZ6AB+JsePgtJXa3xuVFV01V+dHCjlSIyqYeMeiSNI/K9pZAoFysECY9jCtADG7YrLG/0Dz1+e0
eFpHX66ZrU7WVq2nChwBSXPRo/7jfVsKpdwmCEeDJDX8G5fJBMAjzrdp37BM/JKGQ6rsJvrXqHRh
hbUCgg6EyKSDpfEJ7PIoNPtZKRiourJxBt+nw4m/jeqBvW5BNakqaE+E6JFwJmks8UVprMu3Yrq2
fTs5AoRqIdeziBwPELP/Oc0YgM1mSe4+2RdVM/15YYMKfMjd2pcYwcWGSUn2EWW/HMe7qtIZ1HPM
KLEdxvDDngBDzHLKGF257VrE/wbMmaPikuiX8+AoAj8+76/gvtiPyu9p3W3oVWG1lwr3sSt7gMxP
CyU05+emn2U/KN0ML6G/vMrc2rqH9DaY5X4LKTvgIb03z5stezrJhxMbSFPNlAgCQwsOLwS+PCkS
h9aH0+IwYgrN8vb7XwWBGRSWVF/HDB/oP5Mdw9eMBBo0c62iVSHeoawRw3ivux7v3+0fEQtQPF4i
8wgXH/L2dTnWcZ/oc+FCdaqtEI3xZFXwlp14nCHS9BbzhYU0BeD30wp07TasLXqptyCCSxDSKiB9
sQgycOXAKQKXfndHfFoFcR7J2FVi3fuWs3QFCqdiYMiFztWjUWZ9FW1hZCm6HUNO1hvJ7X1d62io
OQXeiuwBRtq0feummWVbULzq8NA2TNt7yYFG8zlUmEJNEYxkWAN01xmcHzhdgkrlVemm01NW/nmZ
e3VTTTjY3yzlDrCktYjigN5zZN7xO4LynMIubxyvJXEh60Uuys6EftU8Hb/12j8r3BtHlqBE6z8s
0BnwkSW0h0qjefo/WzIYun6nIfd8JfDVO3pGd9xKnXVZKjLGyNqiC+pdsF7h9VpYmxWnBVqdEMAR
Ve7WZMYflvMkhioW2VQPT7FxndRzvyLpEkhY8Hrjl0Qhe8XoOdPeUhqJOQAd03NcQYVSOxhDIjeC
vS3UsQmLIHSMY2AgQ7rTHiMutKZs8sfNUGlJLHNG/J8hmSbb5b2j8eQXIa2GXtYiTqk1JyL3bwEm
Sw7n4JGvVPCR8wd48o1ynHC51cB2j61dNPO6z+rdAN8HlnZ8QJ2GFJPXpdOgVQBgOGJfMjZUqpKy
ya83YAES0WHDBogZH2OcDp7ob4RUWW6iwLbHi2eoAjhICqaAU15O7OyCqbHVQxsdEjV1nMlsXxmG
t9DKKNslvFv3xkjkhAA0UV0AT4CO7WrShTmJb9a6oW9ZcbCRbJON9BppMjedEgXkM0xidXzpGC4r
p1JsFqM3tgQmoUuXrPMRQpuaGTE/qJwV/DM8H+rOA/KQ4PRAcK1DwJ9hBAKGBc3TbHPzeF9oZM4h
I2/llDuzEPLvhXwAcTfjDs1n9B7T4UK679yrNetV5s/R1udGh4cIgdgL82WklaWrFRtadjQrcqZb
ES6ck40/MyXBvm7SVnwOXAL5olpxw8Jw6DkKXLm/sdT8DvcvZx0pjXqWA+DmH9zcNwrK2bJfPij8
caR1Uu1KTdf80LlAOfYBAslWWEXIdT/RPehVGkdal4mPqs3K02x/VmbIqext4PH0Crs0Wfv3XeWz
P9FRRs61RiVE9+bOdQwKzX48YyqdxMowPoNcdHa9gPjdKzgqyh70tlOBGAdLRsC2ji9b+y+dqlY4
12w+eb5lld4d6pce/0q8hdMsIHM//3vAdJ9JkrBsnBCI6fLrrb/5K0iSdjHu2/RoNUHJOAZ3wiLw
kID+9AiltYEb8K9z35qQijxl5njkjS9/WfYbLFeY06oP6daMcrHAorlNAopoGsPTtGURA4ApV2ec
QGbgZIg4c+OKxrYcq78GfIfJYb9wQDAm3MTXBAhdgInvPqVeWfMUtA6te1v1NmINTolh81d+5fqJ
1PECqKCjUfj+Um59LjfWger1A/2vBB0QzF4jfIEnw0N0b9Of9CFVBnrKsV6KzIx9qllbPnFqU2mc
0Mn1HsXJK6qKwqzzAu7nhAheLD3mJ+NGzUydnIkeeYOQnK0JlPuU2mxWrUaHZZRCpsdGyA1j5KjJ
rrQ7Bfm+u9w9MSthwu/u/w6rIyS8smUZO/G+IMnOycCtZV1hGmRYx7bemnz4punQrNpvyaLiDgX8
GGbm9ODSt4X310QeMKO5nY5eL+FVFuHkHcKSc37umMMKIwqSqRd2JEjiPbRlyJUejRdOrT81VrDu
xxcbYtXp3VVeIg37+fcfIHfBLI33CBHWstxAFsQONeviW13HCSOsFJQ6SXHkECHe3YPg7Bq8As59
8c2F8QEHJHGJQspwtXhb6O6HiliHkiBDB5p11rMDAgSEe0KoAoCHc5N1AcTlarkVhiX9ybMCG58P
RfhA6vJH+QWWwiVH+YhAZjKgF+ncea2eX61O0VB4zrav8rwjrE7RSniVg6Wd4/ZB8VdcQKs0zCbk
noAFwczwb1LRZ8rOLeKJYLrCDOoHCwYmbR6KyPu1fYwB/Pjq5uQz1Jvd2Bqzv3E1BZ4JbuwEg7MA
wMi/uThINtfIHEoqiQ4co3fWTXowx3YR5v6ArMoAxY5970pG+Egsl1KI10wpmiN34sBmTYHhE8uF
rim4PIahyHg/3rNgIa1C/v8J3PL/H2iiMKT9n0IDFuXSMuhDdi9wcltB8RTnuDFJlPCw2uInWv5N
K6JNiwXC5rFdE26D+5DfyzQk7f/H+YMY8Mm/OqlO70kCFCBnKVIhGnwGxUqxRX+NBl5N79I2+MfG
RxRZ37jSKq6uf4H+jP6p5VgC3iZgO0Jh93uZBFEIf1/8Uv/HmBmCS/FBcLkvSTOeHJ4Y9e+5Q/P+
xZjIOqG+MnqkCw894DWsUczIoBV3ydrbIeC0tReJRIORQLFr4PqaZs2BRvoIJeSH2ELla0Di9s0F
mW1ussLuvVx3vuXrIxfDeHatsSlpmzNj2kl/0bJWVZ+ew1g7nPBrCJxM+thW9YlAuS4Tx3zhACLa
YVgk1pf24f0AP3kH7RrMekh82u/3r4dbO1A6MRyffKsuAz/IgqJOIjK7l//GVgXEt3nml8zxOx21
28CL2J/okOnU+N0MYwT4QeqNOM2lpkLEcKizSm0PFazgfGMOT3ozs6y1oCHYiQUqxktEu+y8+Kw+
ZNdcu6PhiG0Jl41m95uCdVSnIU825Oli74wBRSdnVbXoB8jcFQaLlDBEdiEiwAmalDugkPUxVdgX
cHMizltx0iI9iU3xnZ9+WQyO0Tcl1mDnmlM1OuxGXJRDaYZC/FxuFFIdzCccJbYlqlekxixIFolg
9z0M7XLJQ12YtGW+hn080zOND3mJX2qX9vi3m11K9UZI+QE+WU66ZjxH8/rw+cjRRJncCb4uwNDS
2nxOCqOv3/v0XOD5jBK38VmfUQwMWQBWnQTKRIz3jmbylhHmRtIrgW59cwWR+HcI3/mQCx0Sqj+d
UPnkh8RgGL0r3wfVbZ2Fdarz12B0Ehj3/izkCyXF1kuDP5/oQFeNMYLN7TFU8X50WaaRdCt3iPPg
Q9UTdEiaY0eD22UC49Vt9ekpzWoqZXQYxpeczuZr/2gOpe4fwJlcNj+fUKvReJkf/3jJSBg2Hx0H
9ssfggLfImZS/80qXG/Lcmgtn9e1BJQTYkJIcjRF89S9AvKFnn6oMIkJ2h6LCpRYCNRaB4xy9R1I
+2cLpDXJz1tImVUq/7do9eVhtb0HWVLPTMJ9yIHsqhdbKbQSrD/61I03OfXsnbhsTJi/6l82LPUk
A2MF5ixCz4Ns4XasQpvCm983Tgxz/wfOocohoXwiVxWcdstCAIbwEfNqvV35x5XIMbmS8Gv73kJ2
n3fJhxmxMWaYEVij5ffo1S7T0BvpKShaKFuLYj4O94pVclahmV5gKlg+4CY+dKb7aFFDfYwjpxc4
iTP/tlOs6zr21GreHuD4unFdcMkFipC/K/dh70L05QlK3B1aNQFzsUXXrPwkeVV1jXqWBKSqU2i0
zbMTGtrfQMAx1Sy17/Tm2U4k9urkSIk0nR0eQ2A9/FkNhcW/ea4YVOjcqP1JJdCfS8CQG4tMjJ19
oggs7KOj5fgf6ywNC4N5IVY0kRI38FPSv3ZEnMYUaO8IZFkEBdYEEocb2redOW042AVzaR/TVKSe
/c9TRwgVAzo5720r1rz2U2rbcb4yKiuDrYQoS9tDgUarevFSiZXOfaIwVVO7OBRRorxiMNFD7R5+
2glGWpqaNHPrdrqP36Q0RtqrdxobhRJMzlZt3b6cGiTdZxuCiq8ZgKUFP2I0XjDe0HZL+zz2Ee99
r8foqZp7fOnKRFXJFVamV5fArl0J6ueo1ajkNsbPFAenXzZONBMLE2oIxspRSuB6qlSfujiX7B2U
B2Own5G1pVTcuv0j0c3Y2wQkz7HjKAHG63GIiiyhc8n1HzzvTNoAfGuy0Qs0D6neGP3YREW0FSQq
4xQzKQn45dwfxmTR3Hifwesf0Zx+UR2bgo7EHvccO7XD2AiMhb0XtDiMSRCVOnkk0L9SfWDuKYTY
hA02l9gWzK+F/trk/Rqa29EkzVU4KhyQbPYUtDmD37FyKgZLFlvBVCyO6Y3P27WrRpgnsLGRN4s4
YIbwNFXeCG8E8FkgUB8AxxRMloCf6vAwkE++BNCHGaWw652ZKiqcq0q6w62KwY9yVgFXQhHiAo1d
sKIELonseaGpxQodu71cJFAbZAkIbvshyJDlFQ9ruAB7KR2yaL9mW8p1k1U7dVU1UxU7qZD94n30
sYDeIA5Aq0TQNUqg+Gjamt4O2GRWaHg4XKj5/bqAZZNVB9JwYOBNB6G3sm+Kgrg2T+6mBFUS+z28
1HNtD+NfgrDxSddp16jTubUpIjHfLRYPFU/4Bnofo3sArfIzs1pTHTY1jJ729ebQkCaTMo7Dj/HY
VTs4ai+qQH88XClQSVOUO+THLAiG6mPKjn/OrZkxzyciEPh/gaC+0hGKjllwOM4sEi0TuhOOHjKZ
+y3OutQBnSzc1tcGc7TEizOX+NrrvqupeuAuXiQH14xGpONEZsVdhfBLDXPjgiHigYUwa1uvtiKc
H01GQgENKLw4uKmmjEHo1WsgkAEJybYs2wVqKhSP22LsCtPRy619xxNDyOfGcQQuG2Vk7xD0YGhF
SmjAnO9HyNOnoW2AlMK0eB3Cx7TmM1tQdlG8ibyWuF73t8mD95NRrpKRYdQ5k/9bMzezHF1CUARC
aVb0fiafV5h9zKnjCr1d8u22//gq8K3vHZOH/Rg4dXdEsw49kU6xmKSw1bFMtl4IF1TBR+oQ71VY
b7q3NpmcgR9yJWMiKShGkUdXp0o/bZ8fI1AoPz9az8oPNeDIBM0cehA11ugwXn2ICgjAHAKu/oXl
nDIdGhTxkzJiwk8ZQEAb5iGxCYbsuz7CIWD9hycRGn5NQAxjYxaV3199RMNCq+ynLAeBgkuI2EtN
y6eIHLVIRl3FKP1mOr6oKEehdk+6PgiBQGChFpKGqTTOfMyWjgNzjeGmtMlEOk3QZfwmBMnWVj5d
2v76f9RZqqZdTlJZNiaEpgGhpD9QyEXoNMMuIRTlKFdhFAoiR4QtOr+PtdWY68hrlVxY/N/m1VcU
iiejwzgpi0geCCxhFcbzKwJZNZmz5eupyZuhi+3VNZOdJDQ0SekGTdjYJFy8SfRnudkFtpeZEWUn
MZcQ8KteKLA4XhRkljARXkDOSNKWsgurUTYAUtSaZrBKMze28VWJitm/N+5/lBp0UavkbynVvIFb
8DXAhV032/8reHt2JhHXW46sg/LoqKrMhldBHN+mq0ClaYgSrwQRbUt7/r8AwwR8/MP3Zonyo6D9
DLFs7tHok6vzjpZ+XMdORPPbUT3cvPg7wZ0IaMTkLq5O9Dpg5zheZ8GCzc3IH15PlftA1vpkE8P/
x3Ws7z3MEE3rOzt1H0gSSS454UHpZfbjcFdc+eUERa2DxN2Fr0wNBd3OtqipV2hlWpgSLooZc169
sBv0vuvbY1TOn6+ys8jVSOogUorgZxvoDgVEcrtvpOa7Ok3q5xtnP5+HxaW3wZ40FyadDDt5ol9Q
s4ZAqscftcSgTQARtDySFZNn4k6LhSO/Yyr2bMO+luk7/zjSLH15BWj6wWHrwp6PDGb7VEUVoH0s
RwmvM0oa4J655nol1VCt7CplARKtEjQqwLgpAOqBOzEsgV0nhmH0vY/+Fn92ITG868L293/vB4jK
FPbPrApKEfsvcUX+chFGd/FTHycqy/pSahnaRu8hjyWWdpCRpA2bnMwU/Bp7ihcUuo2hF5S+33K+
uzhkHxZcaM47EG73JwQbVj69zLXf1sQFgS1fwHoAtFLKquaJPsn/L57OxB4Xm2iQiK7N3benm94i
FAMdj/IhxnsGAsGTMM0E9hZN92ZH4MwG5XF1rBX1WknhLW6ykKwlLbD0izL9BjApN0YRixgw+7BZ
Sdim2DT0kQ4AuT8ONGiqsIeDgGclyQq/ePCXZwvWNzvNfMW7tzcSyW1SvvTOz9f6gNM9I71KaKQk
+45vGsP7Jr8LKZnkE1yP5LIiVLJurANaqmKDvt0pIxF68VHzX5SyCNLYFO6i3uKayHTy8V+UTN47
KWoztNdC26/E0+zHaoHZdMarwCp9Qd91LNT10HBpkIkbsTAKosSwRZ6Ed7fglo5R6bl8tvWS524m
6qFaaRLqPLPD6bKHPAweUpQwRJ5kTflht2q3PCHLrkF7EDNNmxblGsIvZt1NkRqzsO+7amSQWa+i
YF+RiF+mGkoJ2EvhpJd57ulJH//BZTETxjMMYdndCGd2ZkRxGfDIvwT6347lRA3Z/IMXy2lT4W/9
Ly5CIlZLsc9/WAXrVkg+2MYjE5qu76A0HRh1WAmmjGZeLCYbewffillWY0qkooetAWPraFXpbpAV
Dzq27gyZKmmYO8crRo0ygX9WJtJpuJKFgVpIt8u+ppiIdv7osTPJDtEFfbkUADVo6n5EWNV+sJpf
fpZcV1j2Xqb1gKCPuXd1biUlwbSMNvVWWwAWKDQgx5eQbAEHC9QaXDDRihrMTKaVWvtG4AReTvzj
aupswvhaSk2AeZndbS2PFlMZCj+h0eeeH8ZGx7uDGXt4zbwO1roqHp6fMV+FZ5oe9nSdZktvvTsi
9yiAyoG7/emHcZwncGHONcU7drpOEGN1T0+zhhe5vCUQpBHrLe15XCB5wa2qKPLCTO3hnehpwdP+
1RaR3O0CjrEPIIIAv+uvQkV8wBvqp13RVuvlC8lAIhSAbYnWjUZoqoU/aN4lGIVX2VrA/BwJRfr3
L1evkBEFkKBOjnzpbw3pEveFOr6l7KiTImua1MYj9gOFs+nzpFHz8aW7YPJao3jwPORVs8SIjoxR
93H+xXIP5zsb9ge4/BYZbhAUYyDyZkXgtgU+JDevv9iU7CF7slh93T302wVFNp+8GGJXrpOsH65t
k9uY8EC6OdGisy143KxyJw9kFgUAurpSTjVIkaCo2LfvmeoEBYdDt1JE9uDFZWfTjzY0K/RRRhkW
TbH/LVKcL2LVZuQgRmMaeg6SGbkXmpZnm+5yBh3pAxOaBfZzZfPQkigkxD2/0kfozAzGIh4XXKVm
v84aM6n9HygMoa77XeUsFT5AqzYtjlmIWlEmQ5IQyNgnPQ0nBN3nFfiU4CUHYOtmkOKCe/DJyZ3S
9CMfDEVm9IfVYMVXou986PlFJAYZkRXFo0NhR1o8XGwtd3iZtDarnZOK+3qP6tREVw3HcsxXRlU0
R5Q+LkdQvRcD91eerSBX/SBb/WM0yUo4Kq0vGCtFhYw0wnigeEKtsLQz1rW+fb8J/RitDcFEpH8Z
xD1a6c2KRpkKiwkxEHa5qOqOnXyKxMxG9VgvMlI7Y2RIjEXPz0i/7ewsSvOBnVogjFv6cWRLNbMM
iOViz35eOBRveypivL7MLN55nz1rP3S7m0MPV+PPLvuFl/mjmZZc+mbUtzEgjvGah9OHtClwXI7R
e1kp7WU4Hrd4bTsccz7fNwsBWoXtc9snwuzjJZalog9pGdNeeM7zIn0DmZpZpUP4r/uFo9GISYV3
rEk55BGAJBKm8FFNbDU9rd3/rhjG8A8PNf1enoEk8YhKiKc/tskEuS0uC1IEY2Tyby3rwrkoMji7
vwvB8Qy2rzYYSaimSPalpG3ecCqiWV+BhIbv53VGRkuvHAtzQ/rm0p0YBgUEwTixl0kaeGieWmQ5
SnRZMj48SRWzTHxiouHl2YrcR9N8KidO6NLyHGeoewCzrcHDQLywmGDu0h6KdBXpw4rxMJwWMxU7
u5wQ6G2QOlBg32kA7hUnEo1nrsFC+Uxly5w6l9RZmws/tbl5XuBBkrd1c84Oimm6jSAxoTsKS7iJ
TZHQbIXq5bgMXl+C9WQbggyCMrAT2PgTlpxkl656g7oCGt2Nhy9NHd/RvqtjFkHesHjSMNOUHjca
4PzbY19icqCv7PKM9wU7ifprLWqLRPZl5yvY1GjjL97Hr0N6j8aMUzHM/+M1+C+g2oO0Dj4B9RuI
lZgI2u8E+06y8CeTaBqujQY1lXTxypRyWm/ynlTxRgGVjhxZtBmLX44rpGfJHOURZsbvogm2E6tA
TPd34FAniOuYay0K/zfy2R8YaR+byU4g78PNzmh/srDmfzl7FATUJOek0470NEGeLBFqX+Ne0thg
qLWqJLbTLpzqr5ENsy3H4F3vfHFgkWoRWLo1SIMArPrb4qYtYKnBnNvqMXBZgIDH8JijP+wVlz9V
M4AinD5ZOQmPcKxNe/RhK7qB5n0eMb8mvO5EPLtveKl6pDz/T9kUvH1oCHwxYZTa660TDor24hsi
85Sk1vBOXYuBJzpf0ue1Rhfn05n0FH7WYlaWV03kmgyyeguxuNy8HDLXZ1OUDO8/VyJb4NLIfMhD
4Ot0Eu0Vgf3hbCMKUKA90aVPxtQmFnwQHsyJcy6P5hOrxSf1hC/XRIDCxB3wy/eNusYendHJglH6
uQWOJuqWAzkdTRcdj4zvkMONXh7VUFZoS6YBUMVWbCicezKjkNlFM5HuUnoS3klhs3LQjCr7eRMU
w2QWMSmV0UA0qDUX07FS+jG+eq7GANrmk1dADJcGMYKBtUt4YYWiinAsvheLmfGfNggZZMZXs4tb
30Z6HuyY1d0clZxcOqj7vN+twCOfUG8wKuHV8SuZNFLtcz+6bKUMqA2Fi236EkZdKtGc9qKBZP6y
+sWxeed3nCGWQ7BmbEZFPKtexfOI8CcRiXFgz0llqPf5QmeGktkzbUX/scXLK6A0UM4qRVkJ8Tx7
TlU2zlCzLiEdmEXlazfTQZf9b884CNEJ8qkrXNqr/OGWUQv12irpkaSuYZ+J+vuOPnH+NHPYedRf
t5TjhIini/aTb4NucWs2rSK/e3M03Fsxh1XCEYtcIKyFhIb0voi04o7ABarWFpm2vZm0r5bzngCe
IXlr4BTJ8DdLDtdkogprNPThQAVUDpT9j9G0s34gbUgzVRtU90gU+vo0eT+gpLVyk/G1E8kM1uTF
MBN+qf4pnZE/oEHIEfLBO99o5GG2HeY4S5qEVMwgEuKzl9dSzSfAtQt6eLYIYBqmqt27YSZgfIEh
tXjpi9g3Jcu0/FYe0VtctcWcMVNVpq0wxTz1KfGkPRTUGhm6M2mrsni0ds6AmQwZxQKb/EYqLdv/
QdRZAHqZhI6cN6zL4pkX1xHLNt/PI8uIAeR7E/AkFRvwZRv2PITBmcBhnM+hvKKGj4A9F9zjSS1p
PMPL8jHHAtxk+K10PI5UDKcX6FjKbirwXEJmlBzNnIZxhEK4ZBLv5v3HA/Utq9I9JlbyPHk7znmf
69Dj9XtxU9mggrUKGQEzCPYmNIV9wbjMqFwvqha6G9t5kCO4AQef8PjA/Cqs0KycRtJcPd8b+gvf
GUCFADXq0WOY0uKp6cptU3owDS5/L98jbRAARBascHhWtSqgy5XNvRO5/RUVnhB9oAA+3Qy78wtP
Kk7BfW42+TrvGD0OzRQQr9zI0RphSjcaNyManNw8uGNT3+xuUwgZPt1Y+tqLSLV/ZAKfC3u84U9F
L85DpHcjEc7Xt3tcOMS+IL8ew+YlfGXwYJr/08gO3rpbTXf7D/afC9IwK4kq4iD2ojCN2VDQ+NMC
KV2g4CtW72H4NAXNyn24Hj8MEMCDKkOQyvyqDb/nqr7ICa/qMjqaECFZyUjGLJ4W5Xjl3SuSCIqF
qYTmq4EqKNgPnX46Df9trEbjPlq7wmzYA6GQlsTI+QzVv/zCDUirXrlSU445V+M3TDGNqKJlpZtc
wuuKr5BclwlJj3zoSUX3n2y/E4VA4S6Ud4r1wDOvFbvxntJ0Nfq6ZtPTXpnb0IW00xzalqDIuVNz
xobU4H72wTclNsYUvmOX1lbdjISUqAy3yp+oXbBQKOnIqm4NTG9LFXLC3nCv3UjI9gFyRXDWpvyL
QRfOO4vF0lCzNCD3/jskhY2Zvaz2+HTEZ56r30UlFjIjguiY0TD/ujfcbXCsc0IgSYXRShMzshJu
AhX5IYRKOp795uZ6s+tMnKx5MRlWnmkk4fKki3RPZVUR7LxjUj8oAE7GyC2/zGjhoHx/XMN3hiON
7pHM5iAlLULvXMCPfeX35yf6eLx3Lelgv3/QUfMbt5xdv6vaSC+6ibj5OP6W6oJBFzD7ZYaucxXr
jchVqZ9t+G0tpD96ny7riqBgIyxkd77F09bQ82m3x4vxlQziujOWaXw+pTgW0Z1uog+5/uT9G7g0
YE2Wq8C6nHUGWwvahJMFGW2njrEQZ2RwJK1J23zEwa8JLAu6VoG92VLCRyLxLZE4FI7ea3u18Wzo
HqEkCnvVmgpSnmpKLNMreZaOQQDbo4/MzVc6PJ1zVDG7OxXJjMmYj52D6xSwLoZb4mycrskrCsxD
skvpZkXWio2DpEnBwy03bn4TKDV/ZN9vxAFhD9aYoCjZND4BwZRfeGi5HRdUKgNcDdHRObicw12m
3x5ss0PjVxdQS9yURK0w8D/WOBBsu42ULMoqh2/cd/dd7RsVOpu7bNXIyy5pszgYM7Uf4YAh1EEt
he69RfHIhopL6Hx98IX2swhWJsvMGQ4bQPRy21hgRIZoNR7b9J61S7p2uRYEHDO7m5jjdY/xcwuO
t7ALwqasEky51VI+trn6SimgDMkpXC2xjTZZz/LRfcFH+eVCLy+1PWuh3EKvjFw4lDYk7CQj4iGN
1/wZo/XL1SWw5cauXCe+/epdOAKRKVrzNxa2+I8jcZoQVAAP8hDJjnjSJOyfOOG7CicAV7te3EVu
BlXDS0D3GoRjRfjqW9yfRZzJFNn/w94HYmXnOC6Om2bnPEDnMVQZeHnUIvGcn2/7NC/5WnuUTlRc
6xXDUsJcEDq6i94R/ZbnZH0YNFzXUikB4wQtA3lVFp9UO0UthPXdVmgn23vs4OTA92ksuimsqCbW
utjGrhfjTVxRSmE9xv+f3591jLaHUgFLDuaJs0TazkKdtfl/Cvv5zrXCGZgo3LXPP+CyIToiUCJG
tj+mneXSthCEwRL3LeSlWrT8dIWnxqMumIGl0WWpo4ZvsdGX85I1mLPIKMHEkHWglpQOtzE9FJA0
VUvB521fxBG0a/TetGoNaNHIU1TlzTMEwAwnDxXH/t6ogVSf8WIC0DAm8UG8i6VJQ1yzPNuZah9V
uaket+TwEb1XptS++gDOP4qiwaOlueJd6y6+F80AUmb4xFBsFrX8Hd1Vld3744EpkT/ElPAZwPBx
lKkN57DjAj1DaKiYHTjEtlKl386ozpA6MX+Rq22sQuQTlMrfruem72PI7FiFmvyYJ3UJ+/4Av4OY
cgncYMv93w2egA3LMdpcMzUoq/bfEoJZUvcodpBJe5zb1fID82Izw/tAVhslQOh2e4v/3LvjwSsX
LlNGQHU202gnOF71pzo6rsUkuFH/O0RkgDO2THOVduGAXuK/5QCtWAHNSYuDe+p0iCi+GLMiC11d
6p2ur3AikTRJEuUl0WJWeoYqWkStheytT/mvvQULLk3Gam0ka3STZIrIzlqtrgrh1AFp1w5QAhfj
x+4Mmmd1+2cc7W5awY00hlBKRY+m3tgylwBrOS63SfLgawfbACKpeAzf4e6io/L0qLHMUeEIiNi9
WEz+18bjH0rz6SLYCD8TEYvSJQ/hXUG65QoH5/Rmsu06ltEhCwm8jkTXQV9qr/VFV1AbQ2ogm/0m
yRwrc0sqbLNdpMDLHABRnYG10apSjT2CxA7PqqJfKrwn3KEetn7LRmOU3XoVVVkdWwB7BKThNLEu
W7WgNHY3fK8q1kwCKvoGLMRacUV5DktyD2t8TbffVXMJM2EyU2sx7VbR2+OeZz3snV+lTzkDunEB
gfBsTt8An04uYDKQ4v+lRCfEnhhWZwGtwnx01Roz1teH3Cvn2GSsclnOwM9t3KYOI1Qwkte6cZuc
eF+BgSNc3OjQ6gVkpxKD5O6Wo5AMFFGMJJt71rK72EvGNvf6K+KCNnY5xPnOoS/MwS8otNbyUWQr
R6tV69hjrQMP/LjHaZwaoC4sowB79AYmZJsXyJcRhwJe5hYyrSu85knopKepqpwcPjUOXrPlMRBw
LJDl7Kd48nkGvbo0imtH+JjASN+jQUj6YIUNh1dmxQkB5xdXAqM0D8vFvrduCI2b54PSE80xnIQD
LArY/qJxZ7/pSdH+EfJyv2su4+Z0vGOtVReSkbgBl4VYPYns6Z+lUXx+feGoRsbHvLyx8McPAGnL
2uujHL1IFrrRpO0Ui8tX8I89VSyYwdtJUx7o31uh9jdA0iF7h7NXF8WFnK0Y7RukUs3w01VUdd1e
f0beI52DOCBSMbhSy4Br5u3NE7ZFUU/PMeP3zxtWxYuvfbGeZHhblQCQezbwYuSjiMxdivTs3N/4
RcaVIVAI3cF7BJPYOLVwFzMImZbaz7r8VlZFo+5w9k6TMx0+18kzGC2R/8HD0mya3iRI3fl1Db/x
5t5h6HbndRico+5RIf8Ub3ibKMbJohlWWP4LFZKJjtSHPJTpgK6H/HAJHqod3BVOTUgLlEIZfKNs
KyWxgYEF8PFR1zQSif/gC7Ma9on0ge948jSkr9E9nzFPuuXmVhe5JYfni8BxtuzjopTf142wkxNj
okxiXvl1IACwdtIVO6uFsAlf0iAV7cLUZHzi6qPEp3KPAO6FK+PlgQnFCBr+cxPSLE0j17xU8VS8
ocfT/tJXJCNlOXQ6DYkD2SJ11uaFTJ2GBMvQpfYTdOHVQ4saWYv3fDswUYPjeF4QVDX4+zYBYPV1
sUaYk2dpkMLrEYz3+6n7mZJowbOedWYzr7buWXOyV7hpyITlfQbyUkzdFlc8K9CaQez2hM635nYp
9rNZhcWRNVPRoRsX41mVceA+eesBqueX0r37i3bG31eM/ekrfeNpFvid6/gP3ClYeQnIlb6JBY3W
YBWOYJNKg7UZJOIIR6chq50YKNauK85nwLdEzNQ8XtiZOe51N1InoLHn8dlM3W0l5ojB5dstQgBP
TVlOoWzRoNGPd67xxWP1HNYGhF+sCeN3dsu6O4HJR4HlWg/DwwZ4TTFPI+EjT16Lt8GXh6mbgQ9o
PEDjc6duUQr6kH99csGF75q07bfgDQT8ibGWc8NDWO2YRUFuJdXgwdwMIK0qFbe/fZi/G1Eps8j4
JsWjaOv1yzqoLsr/yG9TmN7DkmuiCitV/IRciUIR4FFUSA07LqRwvQxYIREUTkWJaaywFYNhg9p5
d9uP7rNXubvByw55UOTCpHWUyiqZt/UWRojHVbv4wMtY6djF4LyNGnXAHAd+90Lg9XD7z5p6HZAS
nopI/xq3SjEOaM640HFxe3gMPEXOgeUv8Lzhu81TGBun00iZSgJvn4FmbBxghb+YVsR7Bo1XSqRY
5cLZeo5v0axchxpRh/bDgbxx86EV8VUZh1s0a1s3THRcN8Udh0zUrTs3ejk109B6C7VEwys5o3Ff
oalEZ0TXv0yJF3PxfoECjrzN46ysSBXKeZadp4XGNFQGHiEvBwFUwsPGbb80UWPZ/knkRJi5ZFoi
ZJhHwEUIYpsG8Y/oaiKREZHNHlDrPU4u3FZPt+LjQD02ouKS6/c2kOoxGBFBDQFoLh3kePrWWoTj
IMM+Kh+hEiYUC9c5HLp4BxS+Z0axsGSzt1uX31Rw+9KMPOp492GIVRu0uEeLNf7X71JhawaGehPu
o1wlfH8U7UMAuffoIJ5ZfSpy0xD7/W/fmfAMh0Zuurty/05JYongvco8Ys9gMNGKDyl0zek4Gs/P
lzGY655GN5QbHjZJ/xUtdNxchQGPhGne40rayt3ZncIyy0iI8Ck6i5nlaFo+Gjp1n9lJ4YgKnaPO
C122pRnwKPackwIZdmlxtUJw3K3rO9DJGMnZKnKaqMnDNz4qDxnaxdWdP/wN70hWOvfoQDofJt4c
HZnHgfd5+Geyc8Cco/PMmLVJsXnSsCCqfdmhkT1bwl/BDo86WK16D2uel7XLTfDRs1BwfChtcjxl
rOC8ssAh8s2eDeCLvIUjzIKIcCH8E+wREHvNFs6P6NEFdHj03Ng1TWYWiM/ihPJjuu8oh3RHi4CP
fyvzjNRqmjGDw+ZoBU5RdLY6hVbZNH0pLsen6HJcHHpsvSqoZ2uDM4Ss52/zQKTG61KkioAaPe47
szaAVo2BIUvbKFqSxXcjYR3jiaQhQUOeyawBFEBQ9tgkc71I85kWT0IgyM7aeh4jTsAh911yR+Kg
jnnHrBOkWBqL5yPIaQ+nlJeHKd+79nEaQvDJKt9T8CW4ToZpnVkrlAyg9Cd7cYpWFhlGgBiqRgUX
d+ZI+OqYbwA6QI+wgjqe8EUfw9HrJKRy3gDYos+Xa80VSO5tDGPKGosIHCgRj08nKSzyHWK3+lup
FMwi+dGUpQD/hzi8Oh9IdryCN5xBt+t6mZuFw00YZwRFuMwSZJa+ZE+VZi9u9UULi4MVHTUmziPc
GbsDSIfJsKpDcLG5pHfdGynDBz+GHzeIFUKijUz7p58zzPEOHIMECtfNIAC3yOhdDc2CSc7wzejs
+F1WpNV2DvTH3S5cgd8bWwEpqJ6vbga1M9uXh4pkXH1+zI7BiO2e1zfoP90sDpCzMFeUOCzGFOIk
Gcdo8R+wplirAyTrt85hkzI6QLvjOZnR9iF1S1UNfshTpGHEEDvUbhCbpF91ptanNUWqmJke4VGV
xmveVrjcHCAiQO0xbhyQCyh4GNkNZeu/Md7z5dfuw5A/bP3e8bak0jm913oOLcer/0d5hIO8uHCA
NbhKPdZQcHbvECHVDHu2FltWjmc5E7/3oHHd3gm5mvKNq6UWtn6zh0sjV7asoGGWkzxnpcfxq6nZ
wnVc90PfKTh+Ei0qmZmqbW30tMAZqAriw4fIF0FIHTSexcXNROH4ND9kktpUr8Myf7uk8oz4I6CF
L8yAVQWR3q+iaKrr6pGVJfd0ft9xge6jxLU5DQNOqiW1WbYfpYoz3p3j6Ms93cdXE3iUUOu2BAc4
8rqLXAlz0qSBgtuTjqn+waZyTzj1Wo3tGde8z3qVAmmHQCX5y8gHHtQIELtpkKoOVx8iW+HKR1Fj
ZDrt7m2R9Wy/GbXyuq03Gvx17c6xaPfzHLxtxRQ9DTIvob4xkCaoKSglTJjKaF0uip3Yd6l+coWK
Q9NuulvgD68kW7WNQwBPL/BWfTNIIfoDL3yQ7ny5CNQB04cnBEzmaA/gotWcnWRuv5W9vF7ZAi1O
fDL3z/uNOafk/raDQQoGT4z9QQ3y+AE94qgv2V3cOLAEAB7wMA9BNH4L2Ul4VPtCZxttS9r9tp9j
B3fxqasT6W0+Xb8AE2eIR94rAN6spBunahRkLx5V0VkvsPSgZJHo9s4nPCRB1MRa+qH+bf/PY0vE
Ns1HzYnBR3+avWxvQcYE3By3dtZkcBoKUHlHKSjWeSInVntMVbmkTLqToVVOU06vezI+FVN7TL28
2mGDTPjUFqeP5jSN6kulS32W+DIbBYYLkUbFBZahdoj7/nole4tY9X+5BANAOedTn/LI8mLj1hsC
LnVayqfmkKk1HI3aHV7u0DANVU1dj3gmeEgOe3oh9mhwXOpp1l/T6M9NUqKE9lsCv1EvCsEIvTsq
MSdxpMh96srjpePW+FcUJkmgXHdY756mZly3rdvUQAtJs0f+Ir/Z+yK3Rz1qsnHeLuc7TyLaDMdY
KgfcYZYIqbbFuCpH2wk12HJIxNveYu0JGhnvArAvgDAWfZc9ME3J6iVSzueNBdlNdPiBOV1UNa+B
va26O0ExiiyFss1+3PhT/k7+M3JAabp+a4aPSVS0K5x3pO1DbLsBRqQR19v+F/WH+1PKTiWHmk09
mchS/fUI4UbbcyvM68vn8/1G+ZvQOTdNejGhJb3v9J3uKh+mKTUQs8+Ns13SDKnwO7b9NKnZSY1h
/AHzLx4T5SqFVo4mQKJD9D568oZGPsNUWeHFz7lhs01WHe2HAmfdKoAiE+Wks5ZA64lW9GvPm9xE
F1BFKGtsLJv/QEa2QO1M/VSQ2XLvP5W5RbhkRx5CgDakESGCYounSznheRxuI3r7SFUyerZt8+LU
CniTJgjE2IRA7Er9yFLQGqNc/gSIPHqXy+UV0aEM41ApXFe9gSU/dSLkXiJYulMjNl0q9XjSd+W5
4KZYzmgaFtyIYYSvwbU8Qs+QLQi4b0K8pRsSNIL+U3mwQX5oF6cIXogpT6IcG8fZX0diOZu5JvG4
R3bk8Mym7yxaC7WWCwNtQbLHHoDvgHhideeTche3JPT2uQrMhsmJvjA/oE39ylMPUv2ZvdKWn9Y9
3DW9ge71DHoGQe3VpCMnq4ZnYuXz6k7rc05bxXOL+XjedBeNiFTftLJDa7n1dq4M1t8jCfWIyGF/
K9AxNsKFNVs+dCzORIgB2usZYI5Ont5uNCjktXtE3oy1AQda61ocCnBetbtAWxYPhmLVuQ93zMos
ICdF78SLOoAPllLX4KdqG0H3jPq6IXyz9Xme1gnlF44+UGyZcoY8IW8a51kCbVhc6KzhzXKQaotb
pIiulInAJkrzDpfe5DqazYSTwqtkO4F/Zz092A3cpmY9AdeycWdaY7/qJUu8hp0uLxqAjzKZbkB+
s43ej/MKS7EmWpXN8D2cIiwJgR0LTjGkwYjYGk3dE16UDdmgNJnVBeOOnIzDz6qiWamoSm6LGeSr
jwKWaI03LLN/3MdboqO/AtrLRL9B07Q7Fusyk5LFHmG+H5SlLd+Rl7foVEl9apdZiohHyf4nmsWM
LdF2s7mEkDSVAW4v87v7P7l+C1H4F2fyTRYNw4wn9NEo4QWpRuJtwWi3Qcbw61Cy6153vbYUMuSZ
TwQ/f7daXRCAa5DYPEfOaNuux6oXrmuE564LpVZdEDPMcZNJPuNUKvpOxMAYxeB0xTkpbcdwuWoj
nsCCG9EV8+RvaBf8EmSwvMad5AYCfqlZ+DWg8u5HIkXTLjM4esTfjVN8/RpZ47FG7x1faVglmYGu
e03M6TXyNoHAkrSGsCeEVH60JyCbFYC4r8L0CoNDVaAVL3NqrOBJA0UsYPCxy5OvzlG76RbHME5V
8e6FEn9I51ZZTweXXgIxvLZH42Xsox2fp4/oZrDZUM/C925VxdWkdViny/zUfx8M0/4PZczgJZXn
s8aL9JVQAwUE/0a5Z0BB9HwMLBpB0+kOhCU7H24JT8eHhEG0cjVRY5ji4jDIIN/qV+MddfJBfWwR
ggoGn9mqwI4hdkxLMAoXEv9bzJdJfk/4n0b5r3+67jK8Va0ueDLypTzoZRyZTlifX/a80q1OK465
3r7RIdLisRXvcKuV/qCACy5oK7S5lG8x7YSSI2wTirgetf/fSVinMco8vLxXhI0jwZ8LdAw32uuS
IrIH+Ld6ck+049LtKWvYm7dSTfdfLdNtPC2l9mGKQ3E80o4DgJX9erK3RuQnWR52baL14REFD1Cb
BdPNO9cMmurgLDFJIgSufHpaTGQSI5lQ9Yx8yHh4cUj5q45ivG1mALazz4eUh/kQycpirvwvGAqi
V+KhlmfnEWksrwrdmWUD4OAfMGCaPJwnoDPG+vb4Q8pPCqOCAbvaAGTguZ+Ffyjws9c/1GgLEqt0
SQlqA4/FXgyBGuSOMc1754aqnTrU3ENmFGyFRD3XS9miwSm5mmnPaQ1VmhPhap36Eq4AfvFVSLMH
6N4Vp19JychFwfZWbAU+hpmoYEuTLY8hgU9Injv3gtK1IW0FbmMwK0rFUDvG0shk1lQ+5vVMrwAf
jxnnAVbJYtMDmgx40e8Sij2XON4yYm+IViaPfhwEWQEJB1RYIIH38a1jD7ip+yTNKD0MuF8I0ld/
Sou0gXg4pjSBqW0VKNhpFWu/Tfjll6fs8sRi7NEzrSpu3IVmUtCdEpnfiW2pqfVgAtLiLwzhiqPQ
ody47AILQPA6xhFQchoTkrMJNGEaZZF+dg4bXHHSm+KNI4VEYr1e+c2Igh93Xk2CMt5owXpjD0OT
49S/YqO35aDdWg0YEVU4eV+vGSROdqn+w+JPZ59x1V3sUHkLcQ0Wl9jtZBWfO76NF0nHQzHxPZsI
w8OZUJ3AUz4AW9twJ7k77gf+RATYFfg9j+0v2AzOCoawaZ1NwVpmqoNXpbDCfMd2aR09kvEJASdn
kRPKKlGCXCeQ/20tko/wqvL/bw0gBAJnNWIv3a3yM/Bk1FBN+hv/2xYEfhH3eT9eeK0bU3kHgSYo
NQeWVthJdtBL47a9FvbhbnAQ/x18/sg9ydAPgzl+NIniQWUSZ/zfoKm1mKnGegJHBlWUODtZdPoV
XTnfBehcSeMy/WsGzX7l0BIiQPVhuUokLSPgV3FwF7qgILu/tcszCozlP2H3qxSeJ58FOFxvLf6a
ByJoTK94OoqXDL5Dz1r7N7+jPUYh+CJ0ZLOL3AAMEFtLL0qJyaMZd2joqHDlmbzoY4VD4DIrI4HU
4riEGKO/K9LKNWc/qzlJI0pcI8kbuzzqOl0LX4EdF422BAsb6BbLX70HKu2PNwFwN9Cr6PR4H+jt
vPDgRyvvVAzSqxO9mohCWr+tVYOLfAh1eFNt/9UT1QuKS1DEj1GQ1NSBijUv3T8+kBw8r6Ss6cRQ
CGa+1H1sDZNE1Gb8Bw55st3DPJuNbAPxISo9XuFfu4kn5sUj7Qdqrqzj28C6skpRBdeDpuApas3J
A7zsnElWPVfXu7wjJ0dxASw0EMWpeH5BPvgr1xGHSlAfvelaHt+dogr/zlJ4W1xOSFZBUjJmE4Tl
hFkaur8B/10FvQOQ860T4RjKIxUvg8N4TTEM6SWoN1+uslb1Qq8Yq3Pu79GAg63JnWCTHh795XE/
oN5qFSPz2OV6SVycpYeRaxPh9ppyA8h58ATrZEB+sVPUAVDPQgMF++rroMe50sxHezj6Kn4HLpQF
yUUgZgFEW8aZ+GAhfBHLcPXLbrOoxQqXtxXXQObgh0fvLaGIRUjpCgq8YdWPtcj+ku8MzidlJ0n5
TNlyeBBl5x1R96DQbD06jZm3OaDrNJBtq4BTYcZ+MGUNSZWQw1h2AnLroMEMheo06a7hGh6lc4Ez
AbhrjSeqFnaSI/N4EAvJSyGZcSibbDVVHxm0wTdRCDSBApYwI5zj5AgItFr496C2x0HHd1lFzZbm
3Q1pl8fiG9YOAYxafBcf8lJyM220Q+3JD5ZUvFQbF0zNQOzXl3aYIItoBBbNDGYTxeXnma50QYsW
PxlVFydU1caQSoKg7gz0ZC+410Ipa7EQL50tHYjYujsObhhjOhL6phVlxBcZ6yH/NdKl9HX6bwcu
oqVuhylOaRhY0fXG8KN6YgbmRIscdV4C5yvchA/Xpx+fQmSwkIfn6qDWcGNT94kZvyukI1k9du15
T5YTZrwHjbzVv852uDcPsN+9AMKia12YeqeD3BZ7FasbL1yhlVInOGPMl/Z3f0QpF56WNYlm1JXc
sqg8ZqgfjALDJERCrKNsh0W8ePLriTIKeQ3tl+0l+ss6hveMEYN0dKtJKFDdcMmWnzmHGH3wbYQy
NfVtkRmnwyxOfkjPCjL2VMJLxKKbeScRK35d+t44D7gS2DjWb34gE88S6vX34W8g/+k9IMPlPpdr
NQW+ACJi6X+xC1XfNcBua9WqGJivkekdPjJUGMOo0BIDG7eYSFsaZwkCvSSSfqT/lcNu7OMf84SZ
vj+OxaLEGF66MrbfCrL5QUSEHHd1zk6rrcv0TBxC66K0koyWn/jsM8onVNmcR7eAKcSTTEYOMBfi
46C311nDreWeMvUuuapWnzbQssCFr3JUnQpFvgP4m5x6h46FQikNaCm0TiBIbW57JrJRlN6U0nop
TSVOzwhuC03w580uLg+HLDGDpPpXB2SvrAzF15JoHCNxP+1fscWjVr+XQzpbM1/r8xuKGDlIy3vg
DeeoNIffDIcNOGiL5FAB/l7EUEBpRV+EotxsyQhwH4tGXVEGhovrUHIJMSOFIB0/2PlprZEb98H5
UqhFb+mvSL10MugxF9b4/M1F9dYK3CuM8xY8gW/LSQRSr2k3+nR8gSbjrRCRfkph2zEhL44FLoz5
gMsKRrVYFSFFI/DhizABoDkLgJLkn8vt0VIZOo9xHgALs/4IOIm19vg3aIpoB1nToBG+oVuvcD9H
IVksY0t3btkMc3kwyiswwGvvzrdTe23pIUrcquzyAjgF7+/r2xs0Xt8Z7FvPJiwFJWLSi9d6GOOV
FgSbbYg0rsWz+IcA9MwQjMhptIuDS6x3B7tAbWxvYZw+TBPUGIAKwuMmGEL9BG9QCADap3sSy7TL
QV+CxFU+qfZv8lamjeAIqLc1RZJjZUO4CPXbJSh201LcYHk4HWTqoK6PBEHleBZlr+7ct5yimkqx
vbNa7OaxctuNE6qXZlvc1caEmFaNv0o1wubx5sp9bOqY47/0x59bHcGDIKyBYPCdeYnw6bpErZXi
Km1kFvNDtntbYxCav/6YZ68MmMNFVkykycNh58J1JciqsDVnq+a3FKw+Qe0h0V7+TCIy2yvJuRJJ
mTd4VOWSgJ6P24Rgk0YZGIdQmt8FHmjQk8hX/e+/kNd7P7j5veytx20zFfHx9XnztzlBqmJrcy+T
sQzk//Za3Dr9rBjyhMCGM9OyDi+ti9Gsdk31ChQuYOPdDgPS8U21YgCGfh8mQkG+utAgSjldv33c
CTXrKLFUFJ12TrrmomGEMQyqWQvSzTHYHa5pNi4jMouTXixIkqzvwuxE56xwJneMrXkY2IBROXDj
l3oy6pRqp5uhs0TjVmTWuPMzg56IZiOAfBWfPgdaV38jkG27Qr1TGJntIkWdRDXcqS/tAlujyEOK
3Itih0Nft2CRzY8MoSxzvMWbPMvicXmzKHh5V5bvMfzFuLbvrVPMEH503JAsviVjxESl7FpqzDWU
yajN6I5UbARrLV11McG/7iLIT8EnxS6Owrnl/H+Wo+cx2wsyGqsp7dPTHFKajTeg+oT7QIVeyKfT
+j/RkBthuE2xGjARtld23oImVdi7UeAwuF/JYhD6Nn3YtuTbh30fI/PDom3twgWKChHTR765AGTQ
BBKgnjVjqUv3KF1E77HJxXkNzlmI52bCE8Gf11XlGxmM4tFnR2xd96tARzM0/98IJNJJN7GTAqt/
Yb7nUSoatemujePcpxP3NKEYQ9iC2pEuPrNMo39rXKgWcq4aZafPVHqmSP/xBFyFRh/D7oF9wAwe
Xg0nAN5ZD5kGrJQ1toEzFBb6C523SLe8Pfo9lvIR+3qfWXMl1YEM4wp8scTtbO40p7Un/sYv++1P
ZdW9k1tnhNtbVE4124qfFlKS9C7A0Vs8A7kAGP8I0QLhhUKAdS7NR84FuLhp5BPnyJO5uIzGTxLV
LsR6aXbBC/83iXnLn5ZhSVQJHei9/puaRcHDIYU6r/4ReX6LET2FNkNISEoFVpQX9YwSxNyWShZO
XQwO7P8Bo4UZVvC+SpSWlWOVLIiqgHEnPs6Uk8XtGq2H294TzA9l0pSGUo5lgFe+WbXXoe4igREL
uFilLSBK3MtQSkJu3ijk9Hwa+uOgSm8puPzXEhJ4E1FLOsFlLT0ZD2jVfBQ5FYAuKm29gPTGDyuC
aMnmEu2TAsCXeTjNk1znyVpDttNA2Zz+4D3L16IECFD2N7WIArWqo289T027jLhXlOx3o5RbQt3r
2LHkpZslL3TdvBkJL0wvgaaAeshJ071OcQPGYH1r2pnYjl4SMaEwx+Me+Lu9kSOO/qLyrcPVlZan
D7J+Dpxkvu21RJq7HZcHpgC4qS77FSRXql02bLlU9NLIzoa8fWf0Hbz5R9Lu5eP4B2HNKBgPogY5
4A0JvcXBq0IE5K5CzVDTgxFnW6hDxckB7o6DIqauQYvDrNBJ13WTXaWIewWfIgJx4EYJOE6Krb4e
Ucsl6HR1gbWrNakGWGbOgQ7u+kiukr8ouKZYcBNtpNWa1Vw7hcAEDoZmgi7H6bY8VzQrNjvNTH3f
1/C2AisYg3EuYvuBKHqQtuztRJw7rwz10EaAt+8qUKPCHIvb0RDh1JPAbe7ESLPkTcfH94qJpLIz
3bXBvo2zf/AukzvmEHCFoNAY+6EjLv+XCVWgy0edA795rSbVXz7isUxEJ0TK1XlV37ry6CzchbTQ
I8EJ2mfi1NGKnEfX9jdX0IpS9q+fC62DbRNMc+mqHkGkhx0jvPcUB6pWcU0Bd+dzRLn/lqua7xpU
Kj0YTvSbi1KSza5Zf27u23eCUvntoBv+eUTz6g4YllDWmpbsi6OTMTS4oTJY7UWAlqF9WBbVEf8Y
3BhMn0Dj+UuT5oB71JfR5tTde6y5oVmpZx3ToOyfd3i1KlAkrxN6z0iyMS9kezE/oMZEbIht1JJq
zoSx8LGGehaECpu+fMtOoZrdHdY4JrlcjrxHMeoJw0X9aF0f80iVdOivrbNwbYdsz0xeqZx8L2tJ
aPVCWV1dAEm+0CGBiwiogWWNv32OEvPnZSFtKvMMEImSRKB1egxBRdFrwEqg5J7WXSgxpHsxz36i
5/I9UJdmP7w3wwaL5wufXRCbM/Un7+J5U3D7sqHcarfNE8qNyQvI80HbQfJEDlpscsSt2ziq09uo
OHYKVGwMXVwXuVG5rZx8KI0103D49e1sPRWsjlJWK12Ol9vQaOKc/I78oEf/XLEzNK9sKvAjDMhB
ADaT76t1zYfYfWcls2mBQ0txNj/qcFc83+E/6C/Ma5B9Optl+jULWmQGVfK4xWPBfYDPFw1prZ5Y
ml/QceHyOpX7weIO+emjpRCgjCac9wyXYyD2gzfrn2vYgt9EJlJC5EZoV/GQqtJio1QhjF16akdf
by9SkNjipVCbR8iejDfO7q518vAhZhtmAnb96yUDyZXWXIviVcu6gXbQdrk61rkqd+ojTkqoe589
+FEZiyz7N8/cD0jH6Ws74HULctVSiO5oH0oJTbuBxC+cKK3zb9UVBBQEYbp2eU1h1TK+kVqWi94U
GVoz2CDoELzrTYaYN9gOU5b3Yq7dHsNWtJSFEuU9SihQMfUx3dY9g7zLHL0mQc4BH9HLSr3roFn7
KLnogLw4vPB71OL80p+2iGR57Ye7Yw1ejWMDVrdyKUqEG2NeC3TyZxqKHXvWWlbYXEQar0+bIee8
VDI5sD56BPb/IHxV1mZA2w8+Nhs0uyemwPqI3oWumBxZN+b34fOV1QMEwc8dUiXHEEXD+YnW6m5/
nxkOzXUFUUz7hXQiJhh9rrKTD8E9gEZmVXqhPRuBuY/eK0ZKA1migpFODxK9RpomNPuRi+aDC4LY
iTF73VuHE+bBROxqd0YbPt8hfuJ5RbFRFRpNmtX/54w4DlIpnyqGyYszv4l7rYIq3hXpRdJse7NF
9vTgrPxTeAB2XLifDGLFh86oNw1yHRHBrfqd67VeGb0+GKfuWc4dh0NVFJQcLYcrHO1j5IaKH4EN
A68oz2WYfynQmHLoLr2F+L96C7cM484vDz2/eY4dU+ktycM8WpAvUNagrLcacHGCy6LH/lp+Lv2H
HDJwUifiOZIi1i1txWs3ExIGBN+UDMSBBgdPMELjYEhibsKvKMSmC440LiHxe1YDtnzSd+cwwmii
wUAf1iIoeOyIzQCko5lFRkLRoTvk3Bi6Ntmu9mAGCyK1/FvL/OpPJ7HAWw8jqHpM5kvwclueatNh
wJMisHw43K38U6qaX8+RIlM6YU1q0i4rT2TZ339zUUxi5iIYGSjrQlti+mxWyHlrp8DUm+FlOj/E
LX7kMO4h096OizTIBJiXWVR4GuPRdiWFKQk2oB4z8MwvPiLewFtfrQgj/VllSRrg3hWXNIfvbPyN
yWaqz7q52rwZR11bjzeccH6Zk6aoEtkNmG8sn+1UdZlEDnYIMLG60LxFvpAbtoUz2o8ih2mxsHj3
FUE3IlCTDufrjJetn8JM9R3VhIKv7o46oEqCH0NpkYvJQ5GzO8PTajBpNFxnt8yQ54baPK2fCbYW
fPMvaQAm6pGti1SbrEELS5TvzuCh/Tebfryvf++HU6K/JuKdBDpFvjqEHyeVfC/Fottg7kPTVQmd
MjpIOAe0kQHDuUpjbV/ACA5TsO7rcSclywJz4/tLfQ4e+DDcG1tppfsMRg/iX84YCU9c/sSk9bWa
a0FcZQKGfQIm08Vp2yQ/oqpDfNz1IvOxLlRnK0fS8T/tFbqtskYkl0QeakRHb05XGmldWkh1cgHR
6VAw9eF0oFG0oHonO6QrEEi2GF7GdT+YYDH25R7SppXw3gsIssX5MZ/Ww6M0Coo84FB0eaFe9oe3
jLJDBudwW7dXjDN7m4ytS8IxrT9oot/0BFM0mpGrFddvxNZshd225rr2MCjIdTJq26oflI+cjvEf
YaGE44bJrvyOlGDRZiYWCqR2jazRpb0v+FO5J8W4O6Q5R4+c/23lUgOUtdSXBbTDXrABsWulGmq7
djL0CFUKazOeq4HvWGdRJ4cFERwjMO+Ul+ruOwZESch8+Dky9WYBJgYsTs21Dwqd6f4LDuhdRoiV
AIMv75sSmH0ASWXH6dwNZL9F5cowB6bdBNz0IeNnf35nC9H2F8WAyiTEM6IPRgCxocHh4C7l8+ta
+XD5jMCgsLKNi7r9uoFc52Uo9THSZQWUjiUpLGciA6q3cH66y6E7NltrS8DvNbZolOrm9m5eJc6c
ENGZ8xItA3VQV22S1L0DHVXEz8CFpr7CSNBumB65EH41GtgyC9aEcU8r2QU6NwrFL4YbeZ7y4tKi
E0tXAE5gnfqavEg3/IhtD9ccL8e03OVFlwoEQ5WSB0m/uNGcyw0pa6JXoFpQjQCyj3MdskWfZpfS
KgctWFQdw4hVTvaUDLSse7qpuUf4nhnu3c/gAUT3x2pNZOhJJ90bR5wKWuGJju3t8GS7ych1s/g9
a55+3wG0K/QHZ5sqDQo9E0Wc3aNI3KTC0ApphJltjpFh2i2DK2B2EjD9QWaLOKKDxLLMkrVPv0RI
qNvl2DP7pQYL0ssgVNrQuAfdja0XMyHFlBTEy+tlfPRDJbuXehSXCrs8Ww8YGw8uQBzFHsUZOWXP
b0GH9YjuBupe8OlfrW+aPdjWd+VVma2T5FK3hZIxqUeoGsHQQbcclKYbgVVIpYwc3kjpPEj98khV
fyteUJPqLAXE6BIz9qt7vgFlyaMBuP0OOIh7UcEau/HJ76VHf8VYy3oTsE2q/fya3eYX4ywTlKfc
W1BIrUdSRzdRTOEZaYofRa7Pnp1b5maXubTKI3ClC64ix4kam2qUr9V/LYJftcJtISgRPkHxNSta
j2vjlOn8vutAKXYVHZE1kld1VsAEICmJvoCGjSC2o4BpPeE+iBh2Ko6mtnCXp0ZA01aH2d3qBVB8
hDxnHw1s0FEnXV3ZLaRRxc5WJI3EifvROXqnBN4YpGDUiRqSGfXCzFRzhCbiWYz1/tk8KqH8TO8U
hKyI8cUZld1xJWVNrHno8WRpkuj9ZckQylMa0w8b64K/yHqHHwh3NFAaIHezT6UNcE0qY5YbWKv+
AU3lNMa+uNa6MpmjQGV8C1FR9IYTVgDT31k3U1UMsfDOC/G4pq11Q6Gd2A3ebeDfmQIsh1/hrFI8
I5lJFevh7WsXdVaUYEPTK9VWBccRGiLkcamE4p4HgH1uGEKaNY1VovzgTsMlf3Xwxpidlm0XASMa
ZGF7Ej8zGmZ7Ve80vMNN4tTiQFaFjkIAGT2aBAva0Tl1yhOaWoU1OfGMkHsg7tDWD+MTWH2eh6Ac
u2rHUQg+PKYgUluRFAR+h0hm5H+1cxuspB4ZwFBAD+x7SstKlIEb8cQ9mGQN1r0OsmtW4RiEUoYS
I0eerX0okVXZ3frnjs0VAiWWX0QkxR4INKbCSJzbqk9kdUYVTUAVwZC/EjiVzwy6K1pdOF/L6CnQ
I5rl8VHofRbe/3HS69Nt2Zs5wAIq7PAtVaWWY8yG+VIOlcfzWWnO5QeCP/0dyBLIk1t/bY0Z0tXE
ylf9Bqq1+wyRUD0oVY3m/PlvswDyllHD99V/951hFgZtm/gBCWaQRlq1+CTLAUlhC4JRVpS1z9+S
qWoLiDpHoKKkhq7be8UUui2H5n9epqfMOQUqgYdEuQzBGzDM4e2LTwoPvesryguqEbESv+VQMw9l
LYjyP/ueT0O1O8YHXRSe+v4MyVEO3QaW1rbSia0OS9fVyOBjuei87S0JRf7SxyG1pbW1WMNNv9mi
Xv3EWf9lJ1M8hdFJvXCDIP91J/jJgXQb+8g1qo++0vGZuRFgOluetRap0HO3pqBHclOT1G1AVm5E
/sQmp9LKeqx0Jp4qOMQVx5CNaasu+IO0d4VTD2D+V+kqd/9eC7PIb3nrvGPgbkPdpSM6Bfq0aZUY
A2j+p72PA7hGo/t/9iCojX+i/lakQEphvaG3Z9P+2OYV8a1bsLGuGmTWmkMdtyf8AwhE9yJvf/yb
9MiE2MXHpythySl7GfEpTqDhDC7lNFBjrXxOyY08AhIG/YyDWhCzSOLvys1SdIV+f64uTJgncD7+
U5/hi/6pXKcMN9GX9GRf9D+3XlqLuk3MpQ0ZfhJQeHMtKlGFx9f5SoSIfsI9n6r3sNBKaAhx3VXM
DkW/lk89NTxSdHuaL20O/1YnNKZXkx6YquMfQNd9hzYIPmc5exr697HGfBBCGdNUGL4gTYuyx4de
NvPAvwHt/OGuGOGeIxEa1AmeieBahqUHF4LGG0IJNkouPcS1uX+2mn28ezJab+wO6z7D3+oI7BVz
Z0//HEwyMm+2Zrb3atBZXfc78PcViLSKj9neH3aQd4gZWkjECWzpteLgMKZvdJpNRRoVR/kc/Bwj
cyaHpqq1HqFtvjvIqKxFS4S1G2ec7o2ZE084XO2/DLgPZkO7mhGK4ugWffdtCXO0IitvMCNcPJbe
ufqqrW0U7zpbIwZIl3pn6atVUW0IEZbcJ3sXl1SvAsgiJE1IEubGl90CYTqhDfVAyKLCoL1tERbh
yewuLIwk+5WH+krMtpUJu3IgKIujiNVm30zmO5GzICPmfiUnIiIZDjQru4NqtAxQw4EZEoSTKkzs
jeJFYH9Beb3yFxxVK0W/L9jxU6Cat5P28DPNgUUHRODlE1Z7CFcJxVp8s0h9hTj2i5gaEUgIcUkl
LxyyhJx7QUFEs+3tjvDxgdpAVJjQRATdUEcOTAd0V4qZwYIrHo6QItjIAbXTBHmzCOfecI4+CTma
Mk4j5x9aC3B0lDTOPvIcGZ7Bu4trWwfOWmRKyl6oJRYSLDOOuQ1iTrTupGExWWJdarJkxpcF5ZWz
E2xRZ22W4lrSXdpgD+iH+uM2lJX1uPxfF9wRGd2xuBfiEaSTXYbFoH0AqjCmRk7aG5gWSvUJW3vl
ZWZj9FjzWQ9nYy9Y8/g3cquMsTkx+15CRv8wHK5Vy5E+a7ml+FVmO6dXf/08uJckiYaV0m2agsuc
3oMzIPMHSX2gmseQpvmIdmAcSsVqSZinp73b43Kgd1B/MRcRU5E1dYO7LFR+gKhNaDmgjw9bzXSG
dJ6NkWwA/nqJhBcKMW/eiK8D3YvbRB7j0opN4X4hj4czqBCEDjhFLaoLAzaFX2oebTap8lPIldor
IEVanShpet4G6RdixSX312K9q6/hek6nsZD8/qlZ30hg6kxRoOs6/8DXYaxNJtRr5zmZha917pEG
zW5gaE6pYlGBKXfoVUsddmraUPO+nVPkzEbYL4AFcLmjdokWQgdGWXxRoVjHzhrvgS7bh4kVdcBh
jWM6kpRBCsdDDg1CXyxM60sYV7ZiCYmmmQhZAcZD5TdrYmlqhIt/1fxHscCoRULqTANBxdDryEzx
Qhv+yFiyHBXvT60IvDgzpQPNnotZpGQvzry/IHEd0sYkeInU+VZ3PoceL5pZjNm8NXxfBiT4NcMw
uPDxEgYr+xnj6bRTkPasaXhw7Ddw285jhN14TexmMTVyByBNfy7q4QxxWXxMVfTGiC/z1Uf/SVtR
1mFJLTyRBJp2LJedAwf+oNWJoLHBrxxN4vpWvcY30DPxw5jHFD4JKimmk6YffeWXwctEZWoRKzlI
hqoL8uslPbW+NWHEmFy2TnYSulrWDk4rKv9pXSAJyElK1blOJjHM1lj95GiJd6vzQKyy7lOukIfa
tFiXSyt79zdFwoFPBqlZrrtedOopV+kV5ZAvroX5ERtRGVLuISk/Q6FLAGPt3mLdRS6h8joPIPKM
Qt7swmdZpDPD2t7GXExHXHlGWhZhWGp6FsvnyIxZPm37FPzRomQE0l9bQDJc+fEGdtZqycizLW5O
V2qZ3NfB3WTIPhldFrxb4bPiJsIVkd9zH+aLBKpSvZq9WODYivYWsMXeTkmoKKEYe/h03seIkWNr
0KoyFssFbky1/aG+AwKjLZKd+amoB9PFzwqkSCWa0tYYUQM+57Z6he3QWWq3grgLcsRZRnqd+dlw
srJVhy6a19ieny2dZkaiui6kdWdixwPu9oLMoausy4uv12XKmA7it+hojjJugwMPT7mQoyat73aw
ZhcixdQWTK6PWNtJgtGlgF92BgX9wtDm3ZTKwsyAu/t6kwVXuGluWJANnx9kSk3crwawKI8fl7IB
l9fm3QCZ2GxQXSqwxhBVIlqh64XqrDEvkbvdMC+ekCMN0EP5Cl8r9f1qMSonZzLdhMjFmVvqbAQ1
7KPTC/ga8Wn8HHk4A25yPRaokDcN5olJHgp47GScyoN17guiN0rxWbftWCPbRRn+47JXbsW3gFt2
wc7az0vENOHRWuvVOtxtBGs1ndTxP3D7dvyQVdT+PMh81j6F5zxoHM6VD6qRa1tJVmHP6+D3TVg5
4gsgCDw1xdsT4NyW7gTmcXOVdTP7NWWzhwrXYLdDeGSE1CkBRD6MZusoL+U4qtVQL7O/5J90RgDm
2N1aYrRRGxiooFGQ0W4EMJBXgkz14sTFpx3/AvVzQwy2v0Yy9PhSzDC9Vm9fHkdvWrHghw9hKjbz
BNM//DQ0nKTpP5JDmRUD0HEvg7oVa5fAjJWaBqw9fJ4IfQeltDqgmqHbL1Hu/hg07X1WUlNDy6PS
KHGy0r7UBK6KYtQffiaMwUdWX/lmgzcOVy1EGXD/K/bimrkbROvOlnESZmoBJCFWv2GSotGrq10Y
hDkO5psp4Er35xYBWguoJxou4kWjy/HsCDzNhkk6lSv4qMIRA5eaaqQyko9iR6kFCDYfduDjohYR
wULTMwfd6caFAYG/VptWEv8IWJkut0vhAgYpBwXxk7pg+CbPpr2N0TuhCrNahBGWY6ZFNDVNqZ+i
LBVBUHc5wUc/JuXr6UNXXpf6sUbrdp4n7vJ4MjJnGEl4Yqdnqn1G1e3DWTpToGR7u//Z1BPsyStE
sMYThL/ZKLurU3Z2ig+MZxFVFiXy5Fde3HJZIkVCXisswlIllDpYp6LavCMdhQ0meiCFLs/sDgmD
ZBGxVk8N8tz7U8hbzjvEQn0Zzc3CVchRfq/IaBEqXt2ifG39zE14gvNhDfoHqMaqldcaPTPMTwaQ
kkUb8kiaFjK8XipF1wc2OxYbn9i6XTAA7JSW/BvKkCJZnl3+KE/ZIvfEVYcrrziuMNc1b0aKzHwH
M5CSsgXIRRaFCsCSM4/cG9EuSW8/1uPZZOcdDEigeV01OBJnkly6nrkz0tiJtsF0JD6ozH2Khuul
ovTNPOcZ65kVJAG8NoM3nUrOmdRxpFMMndwZ0I82BxAWVo5lt9BeEU81MyD2Ps8V9EBUTAs0CE3m
nXw+7p8gVoVdttGjPt/42svfVrTI+++ZK2B6WCehWkKrVvy9yvwSMtuyo8pDK4hnPKnlJMuN+0Rq
BIaj4kwTOzkY5u2Xm45pnsntfYxfvm3h36E/7qxpvbgiyd7zaswAqJ883Ju3PX73P6D3PJMF5fWV
zxhtaPjk0UrrmODer5d9o0GGuZvlZRUkfMAWTsspEOmPqf/RlCg6oy4lrPg55MM4xfCXdCv58zWf
eqWPyO80iUAcznve6F1lusNh3lnWum6gISMolHYKw9DYTeoHqjA6j0MoYYTHSOo9+GXEij/5FVg8
AXLigAHsuFkOpxowsxhYcsu8KBVuxn5P4If/JSLfYTTG69BRFXM7WTHd/JqGIQjr5wei3gPJFf2h
68mpI2REBih1AVHyikMrHJSQYUfad2fguJ09gbA663Kwite1II+GUkQNwxUvEJlRN+W6W1scRFN0
EpEOQA4XoTlEtNTpB6pwFN3bPNvf49Jalo+rGdH/rMgkmV5JD2aVjeCV9WBd1AdCNIJhm3PDPNeQ
vxjYs0xBZVYmYpCf7WcTAt7QvffaIbvJemr9vXJkLdsoaWgyb4DHKI/xVllHax8oFsqEBSn40lsE
RnmEaMKS2+ZvzwyyCrTegFxp+UdXiBumdYarPTjwghtH+VOY4oiETnbXKeWvBs1SPNIl2YlNs+s4
8AIeOd63WHx4mb1eDUEHOiS9zf20aKoDMlWNpbGeYxQmkXTpzN8MU+VFGKnW/TQ9CkpkMaJtx35O
GO159l2SMSY8uD3ZXN9d5vyKrUg9G+AS2hMpseL2PyrJ3tDPzwETxdLPJFSShYqZlbzgxW/XZvVO
bUiLFj9p7Qh3YqWe5Pnk/agJ7BstiKaShDzu1AWwJQP6UnB8dg2ilo4mdJJle+cd8JL+U1o2CToC
MfUVdpl8rMTo1E0opRPy4fUlk6dk/TaUfrbo1tB0AD3N8J+tIEIiU+gvkEOwKte6bab/GB/zN6Zc
lWTlUPhrMbWWL8vzYws06JcEhQSF2n9srWvDofoUNdL+0u/YJfaJR47TEtBeCvXZdpu03zpnhhJG
z7vYId2kzwSWyc57CQQBWrWVugxhXBQcIzfJssjxrM6yTjRRGEb+Ei7bUJdHOPk4dpaYvE0iPUyP
PGiZfvydY9HxYnOygxFNjpBt0NtNACNbpq7rjxFrMF+spiqfJyAQxEKj8gJa8l4+ZGRJJz8tnZDm
VCUZMmRSJzEaKfrfStdx0pZuA6242M4/Tb+4fs9HEXvb5rtQ9LodtNOLZ1n/WUEJWZOHfj6DmVYg
XzPrF14opKnICtZJYsFUZWzkVy9XAxcyV4yhlLcJsaF+JVr+9Plyl30ydhs3SXN6Ud/2De0PMLu8
nYjODNwlH2h4mDTpklDk9lDJBSSIfwC/6eQlzHQulQsbsMfnAK76y94b8cumRc3PUstMHnLzH2CF
s0IABXlKbksugAoS+ON3MbRvvMyPvEIBHKeDdcH9LMpVtY5Yvf+ClH3lBoVH9R3yT+NlDEw5nKIB
lQc91LsBG+3OqUGOFifcPp+CE2N2/sPLuSEtCuW2kg9J4LJE/ZwEGNTjlUmIG0HYoo6ohzreZOVv
RVUx91VYfKMQe+EHWujvsw8J5cD1KyHFfA7k6RagCTVZR2DomlLTZlGXGfRRc6mA0FpAm5dN9xqX
16k/1NUJh2FV4gJ9KyQR2Oa2A28uQ4orCGwRi9D6PiS1j+KtDBkEAYJKIPn9xs5+bRfjgCUNofid
Iixv/3NPueJf+J8hLC1zzsSCA6fx5wXjILhSL/P9HD4ZyyaDur+/ZpfCp/7PXYk/5KMa32Wattqb
k+UVTB/eFeTZDjvmrikqJVgPxccKGWz+j/4K0er9J1nLN368oKXg2phzzfmkYkHq9jgh3reqjNDL
3X0eyTkx/qLWr4CJSg3rBT2QG6/V3lFT6rBKtvE0bjTgqN/qedmaHfOtgxD3w9X5onN5r1dneESx
9gSiCwmuyagqfbuM7G+KiELtyBYVV4yGUhHaxUiONZj22oUYws9YLybddHVAlbnULw/EQIVv34bo
xZxBkhI4Hx6516DmZ67bzLWB1cYcA/1HNbxjyUB3gr9o6o87QoRizshFGx8lSgBtZUi6uq/23sHC
utlW+uPJlSifHYjHTtG2pSwksodAXTBUlxDBm2xWrDXUx6W5FlW6SP+v4WokqxY0X3Ax2mGdg/gg
KhpwXpKifmQEBUIF+rkyF3164uETFz7i0iEdXLdpZ1kTcQ1v7xV/IExCERusAom0HELUpoYr+IXm
v2AIqU6Z5oIV1w2Z/94LN6ddULQEhkHvzVbviAVQjtKmpBbdBH3DDz8Rcmko3IDVsMfF0OKkUWu1
WKrfEV/yVkWWxxuTpA4OzDoE4d82wu+33/Azb2H3nyDNHAEScy9ngopNhebqcD56lbuuQx5htl9u
KlMs5QpzVxoiqEkOruYM73H713i49zGzSkYp6120BpB4w+Gn4kOpmj21lWsv4WjvI8ACCvX5cYW+
+mxlPlU1Oc+LMqENG9XiU5OdqSe0Qaggsj55jLE52I7LeVojjqQMBLZ9GDHZbql9JhErFTRsJQGE
DcZ05hjdEk1JfEOEN1xV7qhAzI6ejWleLqHf0LX94xkWiq2R4r+BinpxPPtc8gWSKwIut88bWV5S
yPY+jNqJLnZCxIgwD21oNLARSNyyQ+fOviUksUmO00m4nPHRYZbh6DMQuB3n8UVgiwhpsaji9pFC
FB+Y+LHByP9OY4AGZsU7XBwDkAuNRKdUChYc5TNg5rOEVfHnF+HMX8XXByvi/5hP1prWtfuqtULC
CI7y8E8ihSd2Q0SY5XxHf05vDPTHzGmZxhO/u03msDL3HXUVcZiY1gfHjHy7deq/jmPb0DSoD8dR
00PNNM2PBxvVCN/iHM1/izHO65k9TtDetrzo+ltSSHZUMJ5ZmXx/Ia1sWmA9DVIs2UHZQgJYz4J1
0kv0ySrgh4SkbOVw+mWEakRXxYN666nt4L1iKqpOtqC6HJRu1YxJwaTmjZBUefKqHCNr93tV1Qrb
7ZQxEizO15gvReyBa23CMV9qzQKUXUfeoiXIGBbCEYRPNKOpDBczPWLgWl9xxsiID/o17oGCdPI8
jIP4gx1PJfyuZJF4FficXwoZk7ofLdJszfxZTSl4cskHaw7RlKOLPSvektjdMTns/tcyaYFxEHAW
ml6xS2TuVFVqZMFZFXzc9mKTvHeMd7plKDk6sgPliE+q5Yw4WIHiNzFVWY5bPFqLiUixwLrEHEpk
5by2h7vMFVur+jCBmWqLg2hiEyegfPLDraMG+CvEwGGYWAxW//m4L8HxTCUqi/1Px2u7Wucqz/Hm
y6up+0lWwG1HP8kfbLiZHbSrDSkoZWX3dSGsS2az4RBdWcZV1eGjBJM8tNybFc9BRsgfSafXTdOr
vyPoaiLNNvVGEEHR7Ivp1S6DeVm4ykmeiBlsL5nEAynrgCiEpmIIrzmzQ3U2d90kuBl8oiISxm/f
X5MYoFxzyC8CzIsKzDqdwj7H0mmsQttt2t6yg2NLytdT1YQVpNX8WiXjXV50VuflV6umlc4DhWsf
uCiJq/uPC9i3DvQx+XW21RGIlnF8Mj55mhHOwsX7svLzNr9InoYkaQivb5tObxRCZpxhlRoMz/Ea
CUUBXTdf5pnbXPifRpYpbPA2SF9i+aS+3SJ06b/a08f4+RDs1oc77KHmGQtYwXphO/IqSpKOTl99
h+1y/HapIRcdUCox+puTq48AF/oStVMQKKE6rIoTGu0KRAXTpwK6gacbAF3bHpzWYq5wq7WoW7Yg
Gimh2ju9crFA5VbmBbr5LdquVEJyaLga1ZkI9GfRqnUH1P+pP3KI1Kb97wVoYKDQQ7rYJAnGg6KE
1YviukI7lQ/C694JO2qFBMpHzD8jf6CGdf/UqNa8t1IxO3KIQ5a82oxleiwHI+fAhX/fvwEtG/GI
0nDzv/XSfWrBx4Xg0FJkJoTkKE9UdbFIJw04bUo/7XYkFTo1L+RrX4139aFrPiG8o9wlEL/SxS3M
tlPtqW926QS0nJNQeyPWPkDpqSwQGdmhxP3BKZCOunThG8MPZswXKzBhiuiuFLyIpm4kt5Jaatq7
8tGx/IBtn0/5mx6zzDv385yQTfzj/tWfZdyoD+SBXTbrjG1/XJvafssGVz21Ar4LHOKkXsUiFRfk
jvj28iq6Ug2+g6wNptdpuEQ9VP96u5kJw7zj9EPp8VLQWx1s6HCK7F6hB3OBIg2wvYmuIEUyUccy
KT0c55XitLz9gZlC6TW+84+wd71d9dY4lylstf3GMGqsw41bjDJBy1LCLpy5gXk9Wh7n2IOVya9K
w9+TN/ofsf5TGchc1367Mvpm/JSSpQTj7pthAbE90clAxgWJo+wptXaiFeEH85/QFSxnE6MW+lmr
13q5PMwH1Bp4O7jYOOWcKB/aFNPnZyJCN57osfbmf6yyKntTRjqoM73nUELBOSp84BAPqZEuXtWi
nBo/2dHppoitmp4GGLjU2ntV2sDXXPi84C224MD5PvOAu2X8X4T6ovTj34G5O/A8zsm1CJGy8oK6
AU9++awYHsIcTJL+KGQPYlwXHYUfpwdpgqwiy/hnTtmgHSBkBNah9JTqw/OGrbDhtqS8WVbsHEl8
68dOTq6ftnp9L8XwpBcOz675m66d3/TPon6E/kaRahHh6RbsYKx1LMr4sWBSyiSVvnF+m8/sTnD/
YnSYQ1jbDWQSqOpK/Eu78bRO3LGULyrupWfSGT6k0Ll43bk0V4YH775SMJfHVmmvZZm552UDSLFW
Kr74WLeYyFT6wkp2icur/cnUltMHuiLLTi5ya9NO3VKGI00QqofHKPXdsAbYs60kVw1NmLoXRV4B
OLSLSFT3Gx5gi+tBABpsLbz9SJJCBrTvBZtFG46c6cAcTfncszlvDHVu6RSVDrScj439j67OLjoE
btZHal1f/7brQFG0BpfC3YSVwFmfxokdclkwKZlwGMwLXQhq0iB4CWan2LJ6WWpHn4xFxRJe1Kvl
6h9uvVBTTiR1KHk427TUQ6XEtxw04DXdOSs0mQf+aW2DjYUCafPRqzqXLoAWj2riqa+y/QemrimO
7tPYioOo5Y6PUvk/h271JWNZeGdO4WHpWL/6c3r1oug6wPi0PaSAvNSht2c4RGKR1c4CWKSlKfzZ
lyO8mUF7gEOWXENtWPXW4MOrdWCro/9LMJ8k1DTrONIJOvzz2b0G2rDEJNWlD3FbqrrIGFUWVm5u
ruCgINVaVDLdD8MX7P8fgB7SPv7vunqmZDbDT1hSC4uQogWr7HHQLNKH0qRZvrh+up1Cc6gFgpZw
jEJN+anj8HtUQcQy9jRG9bl8rD0FtPQ96j+zIt2AkHD8Ir4buu4qxBEj0/G55E5Irpgo0ClWTzzU
esp2DHY6qQZGZwWaLKOTJ1wfLNNnb5OlnMt6wIF7FOTf+HKAl2vYyDMvLqACbAfzNnEzOVjYELuu
98gHDKozYrKH14SScsGfMLk7EbhAVhre5YMnjXC0TOOgxvHscyHOU9R12qTIQfES67WWcomJeVAc
3JeZkWgPtdlgOHDNTjB2oXQKfDbwhEtaKM/Z0NNzCMOUBbCgPFeLBSun1ICkLl8MrKRtBEk5PIr4
rsHGtSJP/GiORhaGDrLYRjcq9LQJghQ9hnvEa1/Pb8kKwgAh0xbiOO7wp044c6YPqJxk8gflWkkE
ezNeLf3McKFsSNGD3h4007RKjR9KPwVF06LZpvJxJXPTroPyipAlesW7BuAItFwLGeiuYDCfROnU
8iqKJwgIt+DsQAeoT+eZF2rzDuf6cH2TTbrRn3V68FGDvCWJFqFQzM1iLSpycpOhufE0MM4N1450
wmiWCnBOleaypXIlaC2wR7IR7kd0RzOgYdPkv9ifmbxIWBD44JwDWtMYKJ773ZjVbe2m34bfLsts
GWqS5k9tjcvKAiwq2hSZKfdWgYXQ2f+AFSpO5/nLWgTG18e19jpf/zJ83L+ehndj9hT1i0yB5qRv
aOaO2zJrvbDmIw+BjAwu3h6eSgGniyeBiaMi4nSDsmPj5GxxzpV+7ureCY0bsN2lnJf7tHizBe7E
OWQsVl9GacjLJsvqo1V0xBio9lFku003wW0RcVXkz7cDZmxC9arU/i+et3jKbfNMczVMaTtHuj5l
1fvq05BTZLklGrBRhqqyd7kHwKgoPYH+RxPgoQ8iuaoIVPkhCHdr1i2nTdSu16cUD4TBn4HqmcnO
WZygRT8tKbL3Pm4CnJTvnguQxcrxrmioc7Mk46I/008Hjpe7PhVfj572x0wUNrd8ruV8idYgPouD
lTJg0xlzD7Ac+CElrQkakaC0OlNY+z97Hmiz/MC0TP1BNukC2A0bGpXB5VakqT/M0vRTVmUblfhJ
U5e2mPlp5TMsJwT/LuJPJLHVnhIMsxlrDcDBtCp7Bv+1pA87yA4VBU9jHKzbA5N09X+XKunprNz3
k5SgPivncUv7rdfS2YleBC1+80M2bU+d497tu6ANic3G1RjrCVxHi2gLhw13WepVslF7OYXNVkrx
OmMyok5PAJUQrGR5nUEi1FQFubJw0lYETYWfQKmmBKh3zdpmwqrEgCTwmRQk44A+5mtWC7xcvKR0
XYk61UKpuisaaF78uSLDve82+Jsvul7WpBqJTQvz1q9ShoL+HGlMfsOQrLxnUtpt5O5D1UPkYvad
I4M23pVEc2I+OZlVqTE4OEckIQeteWL4k88uO7l2eQdDdBz9TVjn9II3Npe5eWETxE7wYaBUfYzB
gh2n4dGmuA6BKhMHzLgcC9eQJqKeXSbxw77sfjUF+rwMIjmnMBbdO1vAnL8066nUSoWkKafUf8UN
6ccvnb5tSEIUfdpXdgSwPhP4epc9dNQ8yoQexpbfw1Wox2s2AQ1Mlci17IV+TPeeje1NlYBvdkCG
kEm1jkwmz3kGDDh9gdmYGqb6F6ApScHSeaoACwA+yP7fumSe3ExpTnyLdUcgqiY8IBdcHRoQDwQO
xv7LAa5NWa3JrflKRTS2P/hNPaORKzB8IjwmTJN4qlZHqB10TfpZhm3MFcY/gXPCxeQ6pSo0Fi++
f9sAQRgz4Pn+/8TIbJvDZuA9ox99gXBUIDhIT0BLKwin79pP8NApqXFe6zW4JnpXztool7kp/uUF
snqF7FBxLJegzMbxiC9gx443ZhQY+WK52F2NpeQ5f1rr0FG2pVBxl+F9SqJJh0OtGfH1ZHksTtPD
OCNiC13tzhY2IhCcbU9TiJAdXybUq9t6noCHn1yAkRR6bBJgcc8oedsgfRxwS3ntpkSmzLavuHHs
4DvNOyI5GOGtNZb0gWFRlSXZwU+kjPNXHMY0b7vlMuPnN4OFQ3hgE8sNSKXW2b3O+XTqQ2blxT2h
NzAlxP2FIV0DjHnsI15BmCl+QLS9B1ifTLyYDU2V3Ol/HUGV50jm4frw4/CLofKsrGgYwHnGtAbC
uH0O85oH6V0JJjzDwLHvG4XqZ9JsU8OwC5yKNMCHlLVJVMDS1CJm3NlINuvgy9IIbC6qRyAFRTKB
2GU6VFz+kjlGLMlLjPoyWMszyuxcxo2RbOidpXVb3BDHHhsOQBnHWnI7MxtTcmIKY3RlE93+PaLh
SWgjaAAVybEZUr9lYZjJveKjUaaeDved0HkzaQ5Ehxu7XHiKRUZ83G+Pb2+QRwQ+APsoqYbmUKTo
g42mW+8iPunTvVZjOrajZDRqYaz1FFnZymJZGun3lxrXJ1wE63//Y5oIdAUru1R1NofBtbJEAqtZ
Ijob8LsaaKNVbbCGSZX2ohXOKrqegYTwXyZPMf/FdQGM/ZDLo/ZzVKgOD7Y0fifeWKsPdTf54qb2
RZ9P3bh/VyladZ9RSoJZNL9721RX4S+i8pGoRAq82kNlg9euxtmq9iaOTeGv/maZFTSOvAhtqeXM
1aP8kZPNdICw5CozyBlx86oMsSjn9wXAYnJ1F5ysJ6mjsQ0MX0HobV9YuGPPxbH2cHKpe1/e4vq3
5ULIj7SvMN51MAQjJl7wFgSdn7xj67E4OXmRxAJ8oR8iYLg5N3qbQerGneiGaQknizOhM/mT0Na1
NgDadEDAO9bfc1zMya1IDCxdxn7PrEMC/Y8T7/ihYlgDErrBVj5NXDcfAo26aZaLwQ+y/jxsj8vR
T+sZBpxLmmwWE92IvZw5ysNA8tK7Inh5AMkT6nx89AAY5cLe1TfsGuIhHP3x66YGmrsEzZncNMCK
C/Ts4gy4GCwckdyJbwfX127nS5FLXLcJ+EOMpbde9gH1OIq62mnyHoWBJjDeyoQuMI3u1/KWqeC7
/w0UAi0vSGq+Do/n0cFCxl/liSvXK0M1enaa9/Re55Q8672y6MU25R/FCzWrmKUYC7Nd96tluRYB
tRLTviBQ6D/7Hz35Ewu8nSJThG50/RH7GGElVcDsLPwZoVuNMoEoSFuQmL2uHpK6ReskxID6ZHtC
pkr8wxEHZWy6mTYcNdVQH4Mz58GtzH7XMfS+70RVL3O+0Votp9XA/aABHNMde7m0IbHoNfK8h7Ga
Vgmk+RS5JDFsPwsCYjS4exgCBkmY2OJQllfxHLkfEw1hYqcVcFa7PgBlBv0ptB8+1qlT44ooaiWm
xhiSVORPCqb9+9rXQSyAFSDxzhd7vYCjR9YPevOa5xn+1NFA00qZZD2lJM8wTLDCiatBR/8hXeHn
sj913Kun8j4JUm5X2kUQEOMxfdp95SVsY2Ta37GFqxQmv2f7H+NFjzCiOyK1PBS738GlwI7ShhC7
NkxEfjzN0CnB3V6pjYzbPHKkxRgdG21Fx0eNYC6yHeS0PJOMh0lowe7WJk1Rp2xEm+fJ21Cn7GC9
0W0QZLtLcuiDoo77l54Wv5TgB9Fj/j8NNsjN/QWQtOZxc8H+zt33JqXwPiWpxdAyUZeSnAk8peV8
MbYhePGb37eOKp/zJrNZ2cAvKU35Mh/hPeXZDhzJQTf4s+T6Kzb4VuxE7RZiep8ZMLrCXw2Dc0qc
uKO2n3sDBjLxe+37uOdigLANt6wrMAYDucgNhCEUIFwdYlmurE93dZ5nNjedl//gMPOmv5nHVDTl
VgLSAoY/pFuZTtyD8f3159STjQO90G/UzBsUhwT6SF75HSgXg5n2Lu+tsWcw3qB38zw9paKed4No
K/6uimzHOCnLNeEellYUbXzDx2Uoh8OQbQ/693Cgcw4zdz3M7BpsfMzgkPkYiCAfn1ELU4jA3LU7
1WoLSWTix+jeV3WUBp7ufaPt7eGSerTsbI5EHyci0XBAA2j+5TypRt05CO8kWDLURWOjspwTzwu1
OKfxaP/7MGK8/06FNzSjd67OV/ozWA9DujSnYJKN3IHtRUYjmltz33BqVu0yYfbDv5GYDgx8RjDe
luwF+cevF479QjP+Cs1pFe7JfzwKKLOoZZFssnrRh0uN5yXGMDjSTbGgEuhT3Fv47rO3Y/GAu6wY
m1EjScIh6tyTtbMrTErxjlmr7P/I7u5i7N8N3xALhJepbV5qCoqk1QxGL+K22rciJZZ/nt5ppzqs
2wTTX8F7JxCiBNSrTk7Bb/p71NsSfrL9NlLia3HwxK6IzKrqg8VSXiKxDksGCbrzUC7VlA7uWmKi
Zejf2mqbM887V5LjikwicCRldZMvx5/j+xGyvQZRrDHUQc+H0IfxZvztDwNeUukx/qhpf2QCzl7z
fC6MLO6FVLQkrRGUgAHJAiQAyxoHLeG6gdWAD5z/RQnIIdMcMMUDE0JsUEfFN6iGUMARemB1srWc
xKB1iUjtVfPkTO586xaP9n+N3VivrMTFoJdZsBMYaEQyNtYX+CHabmrBXg2F8gy8gjqfVi/myfP5
1jPDYwWYzmKKKchKnzFvhj+yupTYBCPXeMOg6ZIswOZ++2NRKGIyMDZcqRgeBSEtUYfmaExw1tgO
WeJa6BPyyBoh5oPfMp3q8Oxq1TbKGFSvaQ91vJUyqqmsZ5kTb04WR/cX2R1895EQhat8nEU+Tone
n+Y3ea3B4tWKPB9WgY9NROeV/VceyIcJGRxRHpOoB7O/A2JLJ0U51LZMsYuJZBJuvcD6G/QvlKHh
kaa1BKWVfvpyoNMIUXcLTT8mpWNdilybLBNRet7ED19+3CV4++5fkGXnIbo+ZaZrNwz8AsvbYt8S
sADKZe+R88izkhcWvKGWtDlAOAyiwOlwCpimd2rjZ/xjJ6LxN1Je0yg12NqpnISEBw6p4m/xxK+P
IbQFw0/fObcZQ4uPBdy8/hjNnd/UY3D0C1+kbr/kQmDXYJQUhIRFWk/3wR1WqokraoqFzl3sVd+p
ZeocHFX6vejqAh20kaxEiERqHzS/A6e9VLH7qc+NmECVNADw9rAdQT6eeI1mK4Z53dYu1gmpYg4D
/Fm68kTiI6d1qqb2OSPw0RbmGY9WasAp8wVtdU1h4JYHMlZu/DO4LNCeRvzo/3jg2lVx7XHeXICY
3pzv9dSWS2G05RJVJKUk0ipS5jhtn3avsFjBaLnKShXB6n0GS4c6Qrw8i4cI1A47ZPD2JR8c8u3T
T6KYdYJaqDZXBYBfnvQhhz1EJJ4fbeKiQPb8/BGiRSGg/mi0LF6EiA2qICTlf8/bk5wuc+hiSIcK
ohGoWQ1yUOQCQORPVjeaTLy+A5HQqz+s5UO224P7k3LGqUQ4P8gHfQo2FoYMSQjvEujp8g+2x2UT
BD49/60LTrzJfIaPkhIm7o1oJ4ie6FSpyF1AUD432Js/Zd4JUeEwpWuL6yQzR1HHZ7ZycjS0ipPv
QxsrVqAdgYTOjMcImBwgx3AqFIbrQ47atIBiCF2MWWKy6Uz0SrQAlh2LK5k3TK1OKjWoVm/TmvPc
f3Qi+jHbDZs4E5a68mpFaXbbjyWRaKD7WKBDLSgeaaX+uTSeZmo2NUr9i8Yekh/+pqVbBsimhJNm
4Mlm7NtPttGV+Thj1+am0/W8Nr0wTEmOELzeVD6YgCdMBSI0cPMzhPAGQJ8Aa2fRsgVJ0nFu2cy/
Y8lWpqv+ojsZF/eEWFwdciQhUFcpMcOFWIhqf9WBUOpWbNgVPS3Dyfieg3FIZ3IjCBu9y6jBka3w
pX7oQhiKPdrqZHs/2A+EoUqH/BNs1r+wnCeIvGjbZ8jTnPuC4EtTeUs2iVEBWbBd/m1xPwfV+P8T
dy9/garY22cHlVXNqO991EsrlwLaciTJqh0WrXDFE6WMw6LECb0mPK9Z2vFqEXOjMKo6Nex0R7kc
rqOnBKI4nA0ceX02yv26DKRPUt0chHUojEdJgUS9crzUNq9PzqEqVagUlYYGlvc6S5j1APiPM2Bj
fvHWHNdSM4GpsEuzsGbRekvHNwhkpf9yXQJuCYgZ8QxuQM9AOScXWuIQ+f53L/YaUJsJYJserk/K
tE64xYHN+4cTA1BOXnQSAUhvY8+z8D12K9jSfNhvXj41AqqSZNtb2HxvERjAmvCp2JylOC2MgYGv
M4Rn/jnOo8k/cg+CHrq/hzH8sDBMjkfi3XAsEEfFr7hLyWuaWGoTuQKaKQnIn8RuHjVKDveF+ElV
8jRHiJrlpDjYxpUdZgngBqoJijxfSmdzCNFQGQrMTtSvX24FHCG6j1KV7SJSo42qcKZJS8r/AGdO
zwUrSMQ6u37We9iqnefiCWwu2OOoTeDAJ1Se7j/LypX7ntlANkcDpSIgV5pZfySSy6qsJv4SA+tx
Pt1Ox8lFpCMA7G/K3/iRMVdlf9c2NSyj9+/H01X9lDniwbzZjNytzLRXfpKIcGljrEmtD5dTzdAA
GBV/5P5xEuhUHpYfpvZP0n6NHx4xg/iEeVEC++W3amjATwIFxTXEoEt5Awt3fi78QMigsROnzofU
iIChzrsAPGtCTJrPU9wEF5JtF0etfFUUy+M3UX89pf1cuLfZvo7nF6N0ZgnXGXrijEyLRY/IA1e2
E4PMtRCj2ZrrFEaeZbUtifXHxqlMhm/0HWf60ZwOj5BpqHR4Y+bruX2qbXl/CmN0uP+Bkxnsuv9d
RJ7p0ppO/4P3Xn0ERIyzrvAXdcvsxcIL2z4KV3ERo7PtpxAdPSLlCzUmE15Dkq0Rqk1rbKcJQ5k6
XL17cfghgEd86WQ+rsd5TDwMjJlxAGSTYBjrdOI849tYtB6lNQmBN0ipNI66I7zPgLX67ekkccnr
u+YkTe+ind3mt7fFsNJwd6lYPXE3XnYEFUHDuWNK+KjIl/0Lm4NmF69GmvLOQuS/yjCukJgxoexz
eax/HfdvTgUXzKVbZib4Dx9koUQ3OzRvxdvMaFAiqlTOU0ZkUw2bVU31KFRDR32xPicl/AaLn7Gb
5gh76LM/OX3/Qg2le5qCwzzxVAsGHTrilZkcMLEGn9IY143+ynTuw2tdBbP3ClosrMyInzrM5jT4
3HEP3w56O6hi4DwXS4i4JZC52v6G46mw3HrWgCgCpSXJuokfYJxZZxhV12paSseSFjsGvVF6NM+Q
Z4w6eLHUfba0I4DGOY0pgg1HBNEKULlYTq3U+B9wLIFKTtfAUPDgS4LlPf/vAX5/lm8Skv3OsA2c
fEApUKKcAHqly0dAlh0PrdnLdE6SSh60Wpm7KnauK6oo6mOV8EPW6wSAKJHiAukiflOIWnQhTJS2
jQ0IXhdsyHzm82iahKSEOfL//gOm0FSGb2itASC/3CEzeXHSJSJcQ+Bx3uX9TzodP92Cjip4VkZ+
Sv3LTGCdMz4EImpCgmzXCC/jQAx3LWhj/FD6G30Mzh5bX19qzRj0hUKTPQpV7ZOUQerJkkpM/Qt6
qoSFmmbCLOc0fGK1nf4xouPOS8YKcy9soXJXQ31/sDSvvJwLGevPhIsS3GqVye7bm/Jy7sMjMA8N
oL7LuHPeWzPWqaaEjPJpYXeLU2aNaQflItB2/cOXU6W0Q1Wm52zIcwhjit//jFCYm5JPic5u7e6F
ij7qw24xgLw6guHNkPuAbf1+tXceAaNoPdRPuov2tjjhy0f+fDsoO5RRRqPGpKDvWyPb48X1HVx9
esfWZyTpv7wiiCd6v6htMJ9mXE8/vaMR7icqfoETIOoW+bI1bhT9YQQtJFDEUuHyvdX24jfz8UoV
Z15wWJYQiLiw+BVkH4y9LljCiCNx9WYjPlVwikgKaQ/T9Q7deS0bLrTdzb2fFkIK7+D2FT4hKHKz
asl17PnxPn1je9MQEjBIST5sw2f3rDQII94vo1mnSP3nCuf4KUR9yQU3k93avpdH9az1k9ENavOI
l31fbeTGDxWzqdFP7lMnaX1hVWa5AjJ/8f6+7OaoKyiretpxxeFvU1yYqG8MQGChS/G/N0nrCSMa
eUq9zcsD1gmbL9PKEVgmuPqLPMKAra6vadEbIGrIIkc4Qasc4PzvLQukt6ZeT/7OsEyBtUXJ5Hro
KAWkFkOYgv6WGgAzuv3/kIX7KyUuR69unKCzxSVwldTXHudNEzKgHQ9/DzYsHW9El/KAe/6wKiml
mNZNI6rKQQxcAX0gqZ+MQml0hU7q528JP+vAGcmFsMmv7fV3knaRN8FxlDiSvxtFt6+s36GcCOrn
1sZd6TqMOFK8nuOOgHvPVq+3zYSioEu45+JGyC4qgSU+b6qltdXxCp7zJoZ/IVxBLqlxcSbpsivc
ezKvNN50/kf7kJAxxYEAX446NtXiTgbEfwDUzlDZOaLlBLuFnpHi/v74ctY74zqnBUQ1d7cGUUod
8+DqmeW07KJK88rsnVFOeHJeB4l5WCU69tQuh6Aswp2nycFHpcmOfdAoSnY/PEMK2ZBTbOOmgzRc
KWWxLt2l3D/Y5pPW/JEuFFjNX3dOhvmalWcFPirgOwX/Xrm0QPGdxzgx3ahQSxXEQyyopKFcZ4Zt
/m5GLlntFfU29oXP3Izkl3epx3B91u3V13OfDmxOF1uMbbfysgqaMB8yUYUWjZXaB2BERM5tY6Nw
tre304rzKJwJunLrZs3dwnfnrOIPfevahJv745SCLyMW02sdU1zD5SoF7MaaPDIt6OS2Xqlo9MXf
oTtgzbyX3qlbI7BfghmN7sEgOUPT8cqf7lRnjhtjLI0loO12LYOoXjeehlyQCp1m6msCTcKJJux/
CboJ4YaT3YpeDz+kryyG67cjmAe87vfLt9yeB4GT6dpq1WLoqILpH2n07tJy04wHJlRM5jtCeWdK
J1rPlKmU29pmzA5q1pv07g08OjyNoyoCIcKysG/lyeSIjna3N35GOpUkDDCgqk1IoFG8T/PHvKA8
rwasMJVGSVOSfhXX8aFcn4rDtOPXuyhD1Wjh0tjtqoj2mXr7J+pJWejDXZ0Yq2qTpd5tgLRXmBWD
epVY1MbOw7MdduV0EtuNEOsnr5V9CvaIIPKQsbLbUCR83FIrqyxi5Nj40yKhjSItYnDU2hTVVAk2
eYvCjhB5sVVUAaThD3fg0tfYXXx2BOMVH8ICU3ZZSiOuSc0De0OAgUeUXADt5LSCWSDVdaeS5NNU
Xj4395JWv7bmz42FjaGKXafOAoFJCdmXC+0l8V6dYCq5Nc8/rtA76z3cLr+Aw1KMoHLi3Vy8ZfxH
gchMFPW27fA10ABBpPShKLQWZgLvSoPUVPdKSCTjvaHuCX7QtdAPbbkdgR1F8R9hfFKcQHWx1W+I
6kjhYUhPZLrQZeYCYq8LbPDtn0bB3wV1K2uSC35sNmbVPsHWNqB9MJMHVoCtkxPeINTUSv6uIrpw
Ko8eWWq1EllOFRpL876d4e1DBELDY6kCfStnZITWdVWaYFipJHmuBMnf5WwaiMBfXJ8UQbfzfQp1
8dxfcRdRSi1513zcs8fhR/i4phsTv+UKfdAUQ7CA428PgJQwb+VXxST2regZKhAWE/9O6/9tHndc
9ZT7m8wyc/41ApTD9z9zjbWeWLCDvCvG2+YLqSKRMpht+NcgHX/2J2Fzdu7DXkmKZzf6Veix5NC3
F7ZAP2wyzJWLAOvoWZZbSPthEmMrNT0GJgS3Hlvfad6b6IUme8xpmkE6yswg9Mr+0UVdVtY4U+SD
HJXIx6BPjLBbPNVi5RKgCfE5eKotFFVecvzuk1UolepnJqGOEkRhxnxAYAOjqi1Ajbv4gQRT2kHF
1bnyG+iwQYbIce2slREvsx1olO56CNw15/F72QjDEm8Uko7FcS3e5JdbbYHD2E0ODXwXD7Po9V38
urIAtBadlQQf9x7RyZfm9+eUG4R7sXvayO8WrvYsWMFaTyoBj11hUs5zHZE1hA1XJPiFgauDO3pi
pb8558nrgISRzybV9hhHd/npnpj+y+oLCqQyvDM3PI5l/3hmi0cQadSkwxp8fhJpeKfErbIurGz9
Hjo/V6R2X/PZ3jLVx+Xb9md7k9A80cgB1pLarAsjrL7TKyAZyp2XqK3ffZi3F1kYLHnpku5UJGwg
8Bfl0dA2zgcLq0tnWCyh+0jVG4+pdfdewgNyTuQLxp1TDN1U6avlYQFgPHKeuIxD6yoWDvv3Uh9i
dnqeEdTMxMcssFoO01/V+LCsFqLsVHxEzkioZD7WEbvcj/gEEPF41HI1OaJ729NcoUjVSxTApDPN
Q2u4gxe7IxtbemQ4xlZmo+Lyvh76qdS98yC6C3wNDRBX0ec2v4zQoPIi7QEwzmzPnOokxmCUcoQQ
ArN9DguL/tR6YB91aEvx27fl3+5HtYAcO+8w8gEYAZO5mgb6I4uALKVJ/yAh3be6rFXn3QsrGJpw
cMPqXU+qZQCrpHWdxi7s8wViWUCPUzhxjJcpQmIyyR0T+1xLu11gif9witEJvSwr/0vQ/MJ74amo
+wsod7jVmgOIimRwKmQnRhGSJHi5LbZCWJ0GonEFP0E/dHWqx6kpTUh0MM1rhyIalPcbCanow77A
27Zmn6mfa7lm/M+m2MuGgT9SOmffsZeIItPKZTMiIXVSVnt+5L6LiKAm9FQvUSQcq0Z2vzhli2v1
YqvqJ+VZGnb4VU9fgG5npLx6hG9tjBSIg0rORLn3drnxSBxX6Kf9Rr06ENkG4qT+e45AlcnvxhWq
YP2MxTOrxOqH54WFJx0eWp86pU9epQ4c4iUvuAHXWcZVpZy4zMofDEdA3ZaCkEgBXkx1fTOaZNFx
uS0MSHdMQVgItfqRvRMiUN+32leuPubC2uqDNGIsVc0Etpuhh3Zk0o7L2XSKdtNdO0ylq7+wPv6q
lFsB5fPaAQNe4zXDB7qwOk43E81bhKyTX30xLO9+xm+RIyq7wIfBeS3At+6mtQsf8BIc8Vz1fx9B
j8BFDeNYpaQLk6L6mNIINrSPj4M0bxR5Z425o80kBkT1IajjK7I709MAsTYUPlXPI1JvRKHpdMlW
lH+5pk5kqc1/6JrAhT0ohpOSsb97jzbwmR6jzS/GtEOar8QKJboS8p83OHErCVb1wCJJc15s1m2J
nM4OtGuUYeKcOGsQToCS7mppP0pvta8BLbpgq8AVirzpTX2M8TG5X7qe4s+oukTtx/wMKu9KSl+/
95ogHPn/cSXI9H1SwwCjKsMyBMEnqm3bqOUT/y/aaaCcIzhZDmnu16NrYJyFnnMkGTvZi+Z9s+xr
uZbDIxQBnSJfS78j1GhTNvk3csHAmXMpOAcuqRJ7x+SoVMpyZacMj8phTnJ+7ijTkMRbHaItrdG4
CuxqBg01rOFvgGODt23pt+hwi7azQ3nFAB4t6AYwuoHu+VszDifzIpllG+uC+kYHyTDXjDOBZWaM
N8meiHwhtwNB8Yizdu4iWoqfaOZeuOi4wpyFGFOfe+2Pr72F8sQFJJjxJp+7l9yyD8/E73zb7oPk
Dt9VqBsLpDhsTO2TkrmlQxAXdIyg4w6/5BKnTlxDAWuczARMkuYFmCXlgJ/Rl0yYbIIfDnhE61Dh
PRRfYdegRG2ltRBHRDyXZTsT4KYfqcciQJcz5VBN/SAZQWA0QvytmOZx/58FVd4zhpUwy9buchjz
oVmKIrs0QMgarT4tRAjw4YpIN4fL4VuoO9pYG89k875rsZtKOOGntmaBPwT0sALaxK9E4S434d81
NipO7tjiaWRQ3cuQGhG1sKxatw4w1rEUDqJq3n0lb3T1oj0qmbx9ca1o6Xynh4CqccwGHvQs1nMQ
HQYHP0Pt61nAx7mkMiPDHYf9sGpPQN+7P/d6WqI0rL69CXb786ZL86GUlg6+ZPO+xwifyDG0AEsN
4t9ExFp0C2aV9SLcASoBCYnZL3l2ZA2CWy32o0JUn2FqGmv9DD2MvJ2OXpc3dnpcYvgnNCz1wp/y
LKhRhHwZko4T2SbPF1iwpEwIZxCiW1yb0WCDwhCw/3hZAMGbxC0kRVHlufPVoYmCR0rKW1S1N+Ma
TsasWboCB0GiFhCmRs+AAL7jdcIJ+qAxroVSr8Cxh3on0B8FLxkyPakM2xp54YWWltfR58Pzwm2y
R9cDczI3o+hE+LUPT71BsGjKAYnH9pbtpj1g9Hu7r49x/HaCEzSNOV5NT6sP2+aY9FwN5e+MKgu7
92jMBNX7olHovVuc8T3aPISjO7d7lFgjlIykitFLl1PzE3jt6YL4+1FHX/Ps6phP/E9XYmbr4krg
dV+yJpIdgxDd2YnXeTK9asKMnPfh6kaUjMX82WkooOK4lfe7LalSu+0HYtdv+8ICrKEcGZm5Mc/z
FgJscj5tA2ci6BtRB6O6Oo429bI9wucbKC7ebcKHjfJEBzGy3GhPpd2u3Ss9TsSnDjqXLfbpa0KR
O7qLmRPVVwCOHqEOmHgjxnVca1aFUdze3s5VOPi5mWrb2cm6WAEhcttuwxQecalg3HPLHPls9HEF
3n0fnsXE/aXUvFMjjqB5X/QQZCkkHJ9djCDgISlKRSz+X4d5rmBjTfzm63zc9CP/3YSZoORZ7zKm
opHEScBCqyyb5MmzyWH2Po3DKLzdPv1ItE0PazMOSE5CSPX3BwiPFGt59UlVMN/3fBrDV+ZksboG
VWfzwpqpH9FICOvjz7utIvDFO4OxhjyzuTYpfvTWPx0Y7wCUOjWkACk/54zDEUbQ+yPVoujR6lWT
ZqIlXiht1/rQoUPSglFs9SA9Bm4aHUsa6xGppUERRhA3OK2JCIWc8J/DrIkKWtIO/NbLOUFdsv7L
4SHVnPMF//WiPrjUr2LBd/j/5OdG+jNcCF5ykNrB8jlberyJkrto98bfbd20PAPw3+h4t+5S1XFm
1KSZjJZgRu8W2Fh8sgN/LvPFoxGlQzcSL1uVOxOcsiwG9RR2dUIuKPDHSO/A120d/AlQoG7btK9s
entR3d4cn4qMgG6xvjRgjHa7+wYXctBDs6CYrpLyFjlInvCAqdAa2a1WWaEbBaAkK1D4cOb2GnGP
SsXeG5jVZmhVyVuT12VrD/LoPDJOOERcxue8c8bUR45lo/qqc8ogKfLHQhG5IdjVe/YJwEpZYrs+
lNj/V654u0U+1lcwF0emNHdn9qyMVa9QnMba135YoLcsE1WG6w8q4QP5k2Ftn5ko3YGdKrUJh59P
uBnE3aPT4jvQ+dfv1FwrHE7r+BTcJWy92EYP8Z4ye3YBSuuik6xafJmwBVyfxwJ4Wq/NmzHassdY
R/xEkDmcFUH/qxf0Ni8UoY3Gmov6qifbHPr1NNir5I9Bp3DRNhRhg4wS6RHHRqvOv8alfDH2bi5L
eP6dBnLe43f7oc/e8eGhUDe1nOwINc6ZLRWL3LAZEKQFFTPP3bW920C6dzyS45Cerag9r3/FuBGY
Gv0pK4psKAgcEGhSECmSvbkoQ2G+g2Fcq9rTCXjeh7uAR15XIU7jjrOTMx1Bwv8bkspl83JXLFiB
TyiQ2dxMoS+GEP9U67130JdMLgEfKEPoggYF8o1FDvU8cE1IyWd4EWM/Tw9nz9BHHg0/s7898a2v
w+AIz/jXG+9ZHOWf8tJfj//tjPLlPbnlyFcqSpb0iKn4CwxpdIpGSTL234rZJEhOgxDYpZdwMo6G
IrwuOEX2yRTAkp3ttRnu5jjVICZZQW7BQYOkjGM1Er39clSR1gDca12+BJ48BfKN9g/QjYEhf6uu
5VSeNjYop7rTeNce6QdL/TnxaSZW7bgwJ1gdJ7WouedsR8bp1kPrzso1RWJyGzq+iBWwtvMt18RE
ZATwh+ylNeVK81+WCiFSNZxuc/xBrwLi05aq/8tdLsw7c0Pdty6wGlLxP/oLgPVE0Mn0+8wIIWmv
O4PW8egEG/n3Aq4ydBQaeCLtr488Ni8TMptv14/avluQLIxPBbJ5gt3lmqoaM/3AsaamfeqrYqDl
sUdHVKQujXL5n9Ux4EhGK6zVwkXVqEUPiXVsNTPAacGc8yChRQQobEtvB70oC6b2pucih7pKpeRi
u2+/3Zq3dLwjK+2pV8f1Y4632oLi3jVQ1a9brUiFBKVhugEJi+taeoitQVLXoQIqV+/83qRhGbPf
1pN7TE7Q9cmJSnL98IYK952+TAx40N3XrrZxXK8yJnvovixv0LBaZo/n3d20Fmf5N/GUKkD1StjY
btkKh1UIb2Zm/ClarR4v09DSMjgxN8w5J7rFUnJmU/PTxiEGgpLt4JvwlmkT+S3N1jrIHIXl1R+f
gWuBJz9svvX+rEt+G885hCMJXfiUBegcutmnLCd6SNiu+7PWR6UIsUqevM9pYj6qojjEmsWNKZXQ
gMfQgGIZpyzmoyk2i+z73Yfpfo5+QdnZyohal8ocBP8lhztLKpdfahRP/XZ7q8PqYndWT4avidEG
aMadHtXZJrKioPIyIVa75ZA9AAUE6+Zs4RarmKxOdgDQe6x6fZXb27aycms4Vp99cTetk5REOviF
f+Fq2aU7mTs3FXYTt+zJ+5WD02oI1F0kybk3X21R2336agg07Tq+pga19Bgppl8tOMB9ccY/BfVI
Ks7CgCmSNDEi8PuCYUb/y3Ohn48cY2umI3ut9zO11BJ1vD8+6qA+pYkGBMV0InbcqKUzr1mXBQl4
wlU9HxvvfBDZwitm7xw+qDTSDSbhSWl0ZEAPnvuCxNDt7v8QLXofvWsmEoMBH0Chy813DVgA28h3
e1jJazUNfDw5ZDceuQVHidOdj2I5Mg4vMIeQtXtY6XxXSCJAC87ChzmrxLB8zWO7Czvkd5d6PPyX
5wm1OueBuSC7o5XPUPbMhMP7lr0lJ9vo/Cc5kMs02XtyWadQHNFf4AxlHLtrP2s4GkQykaBrivD8
x4Il1q/8UpqwPLoflVDy2DpWe062i0wK/SQ8S2BFAu5lttTfMKLszXT2poapgN9YE81hO73jmdNT
juk6ZLESkc5KipCKXhXKoOgjI7bfce3mseBKD6QqnKnTaouJysYh6xiFwKtlHeUE3w9QOa93KTdf
zFbqUcbl3S3Gbr2pq5xlLFQB8A3Qd3YPMFdjX8hYTcr/FnI8JbR7RU5WwR8mynGWotDyoDX+w6el
FbZ8R0G4fxtXINXNy8zJAijbuyh9wrAHFM2QNqJU6phVjpQ6xvT3qabsZmTus+kRczQdXUhoqoXR
WFGdZEJSTMB2GSdCLz40nyNQpJDjLo2xMGN6jZvirl/uCgZ5uJOqqPp2Ia9qb5T+L+/rIJgDfKik
nyM1nWUwgnhEu10NEiNhJcLUJVuATZhINcKTI5ByJPXFrKPgXyxQ3ElMeFCg/MfNSbZAfPqr4Rb9
abYJMKv5LyHx37aGXBJL69MdgGg60YSzBlRtS+MgfmeFITjESILzDle1UMl+JTmrVQeLXhNmOEpU
eQlKz5fp6llVqKv+SCirMstYKrMygd0sKrigqwfapEJf3O/nLs2/nxwGkBp+oh9xfECV5EjU2zWQ
35Lz0tFopulDWipz14EShcVjfmQ3LmI/yBbMgSLvsarwfjxs0posnM61n1c1ar1CvtQX8AAxCmBT
wkOA1AfzxyTTkGuWkW4YyIj3waQoR+TBw3VJ4NbCkqyqH+hchsyWrBpHMXTZsDYqzNKqmsSQXXyR
BcOpSIzqb7S5huEDTd4hlS9bNgUB++6SR2nKJVLUR/JtMGuFCpr+Yea0Ck7ZBdbdPmsqPzKg6AwM
EBRAuIF9vsHGUiUCDi0vtHOMOJ8PtHlA8VULn58ZQQzTaUuoSRggJ/7LnzNi2BsOup1JW0btaMWQ
GAMAn0kzU3g8BpNNXsKdEXE/opb/DMHDbV4fA21WNUl/WCHHVQrkY0CRzOWc2DaZTY5rdqaqJi/+
3MeCBTSNISU6Me0T273hgKGpGPYG4ncUeZbuUmdajQuWL+ZM90BNkqDthWGnQfNyyIkkC4W6RtUf
CvsLZK/WtSp+C+e30zbGQM4FyCPheIOD7Oc25xrlm42d4So9D7N09JdK9NiMYK5uYWGo9V3SXdaA
KAqYLyHrHX1x92rukUXM7nCBJ7t5eyBybh5R9vK6i/2iXIvjxSXynnZZrteRFOvj7IeHa6FbyXza
6B4oGi539NhkrVbiYzyRg/NoCtI8YsxyFXyrY/U7qcV+9oC9SkP+m6fnP6J7YHi2UMEcqv1o6Ivz
ojH/Tu44Z0LlOFFJuewehG9d53h022UzqOiweh9WxmxMZO27CTgzpO2+cG1J6PkcAod7e3D0Ww9K
9tMt/Plewk6taZ/v2U1ap368lohxQaRidCqFrztJMhjXU4Xlbd8HO3uQsjxo2cONj817TFcw/UCe
Rt3KAjK1zGU9NwnUckgJmwGAzTKH5iG5adb6aYOeJf7BTviFVL1mgEyclrDRf1GSN7ms0E7ZaScz
8J5FXADKooc53feLW/kFfuHwsOjSj7NNIuBzTEWQECm+gOkeG+gMnIzQ0Hdx1JjbrZkucwa4203r
9AE8QqP8Xe2kJRLd2alDF5r8TFRg3AGzu2lPcI6vT0ORmK1opQzSUY0ezr4fsnrNY28FShVEx7zs
CVtaRd6a96Q6uQyPMeXMT3HPMWCNV/nT9193zFOicalheSZJVy59auj1O47Vt7OYmcLDvDuh52bo
UrV3W2z2vreow5yONLkrb5ZKDQhyUQHuis3eHI8b7iaEzaZKovRtrhbFhrdqIunTEIvHXeHsB6Qc
GUJXyXCaAYD7lmbQjf+5H3L9wZ838gdaJJBijOeYJU39ZFJvAD08h+bs+rgzFNrBO7H9X5+WizU+
1xWpUA5s2Mx7FGwrwcLBBh3hA1QPA/6Nn24W0DSQEnnoaEMCH+x3nZwPHyLW3fqxWxnI6tTdy4Ka
Hsn3/+9vkztVqlU5Z/K8ngaMbGSh0nDhoKeDMsH77u1Vvc0TaVfnl6rCDMZhO9bVjZLNwBRzFtdx
ztHz52SmaeaWW10HPeV+LkDVnJrW3L/FmGdR5aErh4LHjXxwXFpx8uuYnBFSOVLCviqLD2IlpjYs
CsY0kTI/uqUAcXGuSLzBD2GFvZ+8EKnKs0H17JDsx1fWmhcluHUR8djWy0J9feARaREW25aNRIpj
mLnuCj5Qi/A/oM8CW1fIQwwgxAILUk3zQ9hHDPBhP95OIJj940P6Zoa2HH2ZsRM/evbA63XCELys
niRE3T0XCvzk+Jq9Nmc0n/kSf7SGCMKIB2OSuhmPJd1horjKm2mIIhV/B9Ojit3E58soE/xK3eii
Z6RLDWnEsPJtEdqhOJMG88uEONTVwE1NvmCI+6aaPlIc81UPndikBWxDTN7stj94HiUuzrxg18lt
ZAIw5LRNhkzUlKoyN8xn4GqDOuuPS1VUUlDsJon0M3/dBeqGJHQAfOoIIKO0ZJIEe4GiY0s43Vma
Yg0HWXmKwsJMwNdvcJkZavq7WBRSh1oxS6Cw2zXreKewlgqk1d6PlE310cq23yYqBm/ds5k9UCCG
L7PG58cx/OENz04YZUkIP9/XyDnlwjMyI6Sqm5C8W7ORPH/WGx+wJvku3Wz3WuLET9eF0gZNf6kS
bQcJJbHrIYbAFK+iDtjvuiH58nENa+TM77a/b0E2x/AlKnUvhpUP4L6KrKOgIpYexeLQPAqaaL0Y
DsQE6U4lgq/wIqzvuT7S6TwUM+RCsW2vIL/5FxcDL6AY50uvuxVGNtGkuFterzywzFP65uSunHYy
WL3i+SC5FSyjOxQulLlDNj1HgDjAktRvX5cl6Bjvk6j4ScFoLxpX+IDGuXcLTfAUivOWW5/pL5nM
UWB/sEq1vrC0MI6dFffGlVb25XDcLtPnvfa5m829SAKEW5f9m4X2Pk0nfHGT53cDckaWlc92MsBl
0GsCQiprv8Stb/inivYQrb+rcxGSS8gDdKnyVl/xB10pLL79F273QDwzid59klYT+pd9lG4efjcf
JnfoRv69GE4z3WKSBQYyDtQUIMRRjN3/6WvORMhGAYROxdxadQiKLBhQqQlx+GWH3yt9rHGQKK2p
neQuni8La0BZHwZT0W38bCPX2y3HIHDIxXshgJvoZI7j1ol4Jqjh0HOrgOia8VtFFcon+SElghHl
eDl6OgbBRbr8ozINkjsO438B9R700XPMnfcmy7+73xQRzGKaNTp92K2uZgZyFGDPxkLGyT0HFhvd
kVMSBKo+2w627WNtBe4p+VPwwmh181IvHFoC83T1Iujcd6wptRFajBtSL/UZ/TLK4zBwcDfH6cor
53hyyNjolD1+OEIhBaRQC8sfvjvYBpGiLVXmvqZNXs9jeEgi6wM0KGJ+OXGuiuA8DC3H158pPSaf
cKHYW2LtsrKqAZk1iQfruygIM3GQjBqFpSZfnfH3gg0DWoNA5y7V2ln5PG5wzpOHNGCJCsGNrwDM
cUtJsM1c22avMpcKo9zXfeAaA30j0gH8OOYBPhHiHGOeiW6C9gMFv7ORaLWKpTP9T3jJAMiPq1Zf
3fijgz5wrc31fFxQ+f/D/ChUwv2YgXrJCs6g7o8UUn73L6s6j1JCuOYJgJ8nr4WHiu+WbXwLLQW2
XfmUqX14bYKR6MSiBKS/dC3hfTlduxgVEX4z9x9cZKbEMyY3TFPtbAiGpj2tDohNjwSUfsLnONg9
zWzizVZcmG1W8iGSNejQMDGwe85uuotZX4BA1Oi0iZnEsAgWgjfZ2I1SwSlNlI4eHim1JVUZLdXd
H880INDssu/R9N5avoKo+/exDC/V1asG9RXFREVX4FGWnHAUHvzZ555EAX2pFSKpFe8MXrVhJj26
61N8D8CqOeB+hlDh7hbDZHRDFiT4UoVb6n0DMI6qnl40kJpwgsPjJqbyBSc1GQdB2r19BlgjouTC
C0lPzShPIUX+oZPQF0wEp6vHDy6yOeUrqiOFMBe6VPS7k4Xq4N2UvAOmf6iyyM2zPDGHX9Nzu8fH
B8Su8K3trolZWNHnY+u8oSunk8AQAFN00Hyp5ekuI82uoxG3HKhRRZbs2yl6OsRV/vGJis4Hm+re
UAowkJxp+sObfa6BM1g1xX6GLTkUnq5LO3QG9WJICA0O+QaAKiwRVWh+2qp5M26AltVzlAJD0C5v
PN1AaX9NId21n4cLkD9a2UPPSuFSKQ5W6iZoZlxZf/EdLr2LAlj501RawnTBlzUqRzTUitTjILIu
lgS9jsV6FA8VYkxMvIhzGS1stvjfHbjHfkEqIWPoGA9TEtnzYZzazcsC9ijH1j3/5Q+WcGffklbp
E/ZfgOf3S0zIBoY1K+dU75MmNSYxwO1mWobDW3CHV6X0ymPfPEMQvTvDMvnF58zGpCChKcLT58bv
+I7Zc4rgpFOvXgnkjHNbpVJPB0Jydp3qd9I0h4HwI7cFYU2dFKG5T4pdJ8IL/E3LliGBDFLhfrgM
gvBKObf/9OwdObJgQ+zCobO7+3uz+uLe7GxTkdWCijaMHKonPf00shIn3J9IJVU/mKkbKI63xiAR
anPrAQyGIDLpNm8c7fRSOPhX23AyF1ijHX3iCumDIXY1rD5ONEWjZ1q59M1EU3T2rwJrayVBimNj
ZqbFrDJITOtseR1W+dtUxlEYzD3nCuZhB4is6n3FX0HyOuhxKVKi7MmpnUhIl3JyAyhgwqE3uu6i
/GdgqPxpFGUSfz92Ydkc6Xv0vVaOB9kpX+llF8E3+fvaGGkTT9Qt/CCcb425nRPI44vfMKcXWS3O
1CXNLCEtmgjFbTIsxEPk7nPWhpU3DABn1DwWIfFy/59WycXKc9o3yDsCN1d/DvW2tk8jOPNhbj9p
Xghlc9B/v4hcDbzMHJapDkgB+o6Akt+sG9nnouE6LfmAR71pp+fx50tWkxoFy5JUyGrBEXYDTdJO
twwVXl+8BXp/GLY6mJ9gFwNPF1EIh1I/UUz0jfNEg/h20Q2yS9QFCOaHIEcRCaD+pcdaHxS45kED
EwjEcWu/NR9GWsIYMnyJUg91hJ/ZY1Kk0HhprPH9gjY1DHneaY4vuKnJT7IGluwxmMzEoSMH+9fJ
EqvVvugK6BpWbhVcKPgpNb7vmVFT0F1r+cCZq8NGlIU584LHeGvOLyJnDFS9jLQuwf1sBNdJ6UAv
WMx1+Jnsygo6jzdjJ6t3FBthIgYtyAQK3hMkaXjCv8ON5ZEqV/R3gQqRE+yVAynWZ9734OtM3MBy
yx4dwc3NHdwwWyRN++IMM8wWO/azUTb+xLi3LaO9ISFMt56ltIx1aQ4r+NELk8JTD+QY3SnnqInO
IGy2ixOEZs7UXj9lgovTg76TRGhimsyzpK4AC/l+xhtMIl4kmYTuaqjaQ52jiE/PIUl6rnPqamHQ
Mupi6iHtOk4WVA1UYkfUrWxdH/NG6Rkyjjxgyzznmx7JcU9tB4gukvuCKWC7IkQGyVpXmNPddaFu
v4atHsEQHMPMeiTDUjwkuUlZ1kBRdh+oGfwSCG9/qgZ6lXZBi73DW25Z4FqEyGQp2zjtIxzCwKc4
yQw+TsQA3hsZUYvBnQW2nQ3iMTvnYQsJyTW+RG+qN5ydRk7M/5o451JDF1p5dwVP48fSCtx57A0U
7l27JdIyXK+LervQjBpLiBBk1sRJOei8vlzeNTq6F5jPcdbN33OGE6ZiCKTtw5aXmYRdCISGbjBO
sEdsmognEb87u8vNvMxldzG444uIJ808Pt1JWYuOaptJ3YWo7Ta0Cl/yDke44hpvynJtgka523Ma
6QejHgAa1diQw+xLV8RxkczWYGgbcL11J4sYTGTQ4IGcA3SaW/mzXlKxJMvaxpKyr34+P4ZtCkyr
FcsXTiE+/sLm58YyrOMNXIhCWY7QS8f1WaPu6jz7RQwBG311Wedw/R8BLXOCLzeNlIDuiYR40DKs
MEdnAVSITtkRzXHOOdx7TmQdY0dlbw7W9wd70wpSd39DlRDN8UwIoKAEk7Tkrof799L6XKRSV3Re
ydAAO7Fso9/evEqnveEdU2QQlEXTHE+V6/KlCZpc4IL9yhK826PlKT0PKVHdV42L5K/SZBAnL974
1gaPDHI09+yFFWJKnkribtqbZ5T04Lod3HRzNDkdFCBSWtKt9ZuyEUQNJcjbNWpZ6o/xtrzMTddK
0doLGI80rgwAfNDCKCkPqfqO/pCcyyui9VM64lL5JjH722TFeBy+KJS9MRj1ryg6+MRDQnss9fDP
iDJPWryU94vzJDacBVURhodn5u68Qm/hSErDNaxaB9NL+jD/E2+2pdDlTrtbhuJmtAmHk0vscymK
xl/J/mmBXoh+HhnzUM4EscD3iGnNt9WxIYtpLI5gIH8DIS63ojs9sqUFbRcCtTPf5VXRb7p8Chcs
f+I0KH+/44vVz1bsQ8NhyochSTpcuJlQHS+8GuY87yuVGKt/N9HXRVk08YC3R54huAsVmGACwIyY
PglXOTTzrC6Sz0Oa1Id2g+ZmAOB9aTPr6ouwf+eLQem1zGrkwtvAg9cXw71pa+n2MmU0lHsMbE5H
v3K/qj9ka2T5EHEYINJDHw+Nwhe136C2M7lmy8smXCsEEsJrS756/WgHlfxe5BfijTpvXdfVAIHW
kvmBSikvW+SJDDr/mTsc1LUVa+uj+lq8/xk8Od4973woUegYstryssCenbxv/l3xdxrgGN7PcNXa
2oS9ITceVaJhmkYQsbfgL+IcmTMkqNj9hmU3O9kI2xvsUsYG4jcsZjQ4zI35JsZcEm9xBWV/HUqQ
CIp9MP2Si0zJQPRHgeHB7Sq+dzOBSjASx+GO+6WoAU15GQFUH6om8nx8UwRe/msIEfvHp53KNnf+
jH3wxw2lYN1bAFwLWBytGDa3NrVK3ah0qvAOFvb+VyitRY36yjQQMJcyekbClR77itnrOI1NL76E
JWICgkO9m1PizckiCsiF4HlzIXac4vcq+j2m7YZ2iS1fr/m9K/+TUDATmnSN9a8uaLSpYddOKJWx
vgNLbovAw1aDaBMgo14ZxWIKLbsyOpB5xc93JMbjjphQkrzGXxblm3NGvnojAli+Fi7iqqmOu3WV
UAARcdRL8aeAL6ukrkrBQEzOjo4VBXNd+AIegYONldQk//o3nwR1x3nT9ohS8qHo8O4/y1bh0GbS
3rQJJ6NNAS+kMOSbtwUayLtP8m6P7KDC+OLe4SoJ9/iuqsJHbazuAnsc+wYqUmRiMynUSfjVhTcR
HW+LJtibCq+BVqGx2gDXJgTqFeD+YBlLNd/AMD+H4e1szgzg0jCmFMFXy25VTSGvH7p3uj2D0kTy
oSVUEiIeTLQWg3QuXoftXPqNzkRBfM2dQ5psjcjmthP6wwxIvHrrTVcZAJmB7H7GlqrHZXGuOYYT
mPuANLYPB1MtA4CIx2mOnRkHMEPJVj/XiWVbxGIqaWWgLQIvmT+ykke0kdc6yT+rF0OTc6YuRvTj
/9WshaoDivDlKwK+y0YXH+uWqi894qDRg4XqFYYktvOexid0p+vH508OCFG/WcYmHdjWNJI5WFzw
/yypTopXhYw3s4uviy0DOWNqL4H51LBtf+Xe+i7Sivnsp1kT7jah/gHxCm/JzaDncXtXUzSVGqH4
6QBXFLpPs+LxVvr+TpVq7DYsMC3Ry6HUG4WtsWEuE6mHZZnKTaoY1Uh2It9aHHKlnLuhhZGDCZ3X
YguMYAo4pVTxt2Vuhi5RM72jAtnIUjj/NQmd38k5tGL4rXo9SJXpWr1EMFO6bE8qH7U7ReLlY2cJ
l6qkjvwK4CMns5HJjyPdwaj1M3KgYlcBLqJP1nNTxEz6d/GHBNJm3kxw4bjvDB5tMTRHVT9Ek+fb
p3ra8cUTKd2tVMrDeGjBrGGTu+6gAnDQspfwcgZRx1oMaBrSxU5jjG7dETvm22YdV2JH08g4Glxv
/uFpLJfnXts7tvI8Q7E5Yys4HZbvGDiGeFUXDcGOMYExUeSIx4yGxmiFezLvw563ouIw6raRqXa6
/udRKxE9EUceeGwHcvHyRYHh5XmgTxWm7Vp66wKRi+WnOwDyhla1UemykxZLufQXnU8Oz+a2Cupv
uYcNK1zUOIaYtr662NdBjI3olNUu9o4j0Ucr9bVAcsBOfCig/9gjKL06plj+k6Th78S8iahnLsW5
pv9fnAqRzyd0Z87YM7GsgelK7aHa1rPK/zZczHdF3hKTdb27hAZcnakrWGWuHxiL1Dgnv3C1ZNn5
uXjt55DjyVPPH4LePpee+AHOBd42F9BJmA7b1THTlBOgw55xOIGiSb9VgmjWr+ZsGuoMJz/gbU69
eomF4aLvmMAKVdj6iubOxyOB4jeVfEI4oCbXK90YX3eQ1x9IWYpMPjtUu3VEm6q4cdc3bmEtiKBP
ysUIQWUl21KF69WqG6Kbd9d2T5j61Lv6hQNqTuBhWfZWa0/YfA1XuKBeFHY6W3UMMeaEEbKD0uee
9ZkhaPPJ4TvsNfyMaTA8EnFXbkMXJhDxhQI9gbj7M6HLrL2D4nbPzolIuals4PoyPmEuO9lgZEDW
aBzrpv6O7LTIjermlXFZbI2TCtJ3eYFrFPa2pulon7Gf1Mnpf4MrZ8wOfMXPHieJxzAS23nCqgC2
eCb1GTymhTstGH6drv0OnAhsC2IwAXulxcjR15RgrwM+k47cn7zBXMDOjgyui66cgrnlcJm9hlNo
bttt+CUJ1UpZgdT3722lYrXU1zcKOQ82T/fF7atmue8qIK/Sx3ZAh6AO4DBpjbDpC6OyZvks8IOS
QFJTzdHJ9bxBGFdyQyAwGsQa7et9VJzKkiUstZfXfeJoSUPv0BGyXUdA+bKsuVOr2u4dmbDRSooh
+whynq4bQLxMwYBOhnv+iI+z7PMFGVHSc6Gb+9NaOH3OGRv+boIKM2ZxxoHLcVJPbNbUAUgsSR0O
P9lge4jQE9gYnGHIKZmzFUtiNYCeoq0f4Vgo7wi9Sw8svmqL3gQ98o4ve1mB4FY492u/E8aJFZJn
gGQrdJL4L3K2y8FxNkgawlr7OPDMYnyaNk4YaRAVfgtne1iqsjxgZL4YpcO8LimDXSkmUj0qEINg
wXHHTbMaoMO39tP/3Zkpdf8yFiWVYHFp06q/k1RXsi2HYmWd5kwJwTpZMVvAakWkFfj3fd/CGs2b
tUWK2s90i178/bqq6UW/xVkbPh3RGpqwfQuBpwqzo21KTnhgdH+1UeTxEEYAc+YD/+Pg/xdGe0zO
nS6qYBe+YLOCjIY2uOg+xKcp/1ZuKw2KrS9iGxbh8rbWGOZz9sspBfAE1sif+jm4Tcs/AbxJzuvp
S2bbFcSg1NPVkEYZayMdYJY3VSee25txUIuq/0er27rbnSJYLUG+fy8HNQpQOM70wrpcaOu0hroi
jGsbUS43J3QPIBhKDt79wqZk7UAl5TIi8zJpFUdYDxCubaV1t4mzMNWlc9hTuV7zzpAJEjC8sD6Q
myBT8eBrQO2U3w/kqTttWmwOPUAayUgWxpWDvLSjW71DQd2jqcFzJzHkQdcv6wJEV+nxMFFtSMXh
Up3iM4AkjfZcuk7B2sgXb0UQsQhv1/X+ZXEHhRArltmFZb9i0fl+7JlkvEty2JSmhavI/H3DW8ag
AO3T/rb3Q1vaij//YaKB9s70VuM29OV2ZjBctbMcWCxTkl4F7TKPykathOioGqMihGQ0g1/q93HH
fQlZd8EGIRFDU9opTEOrfmUgikCe4AswEvb2Mm5VVvdx1FoIyfveit7xQw5H/5u4AzkolOuxVhXj
E3wVzl9REEwfuYDgJkn4wHhoIAbde2uEAcW8qwdKqsMZbvjgdGt+AYmcLi2XxCzcdzZ3URRgdAoF
ibIfSO24rAff/VKf2fJQMTCKrnwoIUGvffNwD8vYlyhrg7A9EE7Fd2w5m4ln/r539DMMF6XptYuq
9D3E7kSrWUIkrmb3yR/gX34jIntgPeJey2Adg7SQMAsJ/Tn/VRp4wm04BDO8hLmmbtfLF/ycDnFj
DV3xFotn+ldRzQGGF7WJF/N7lQ9LoOH94eabLYDDy32b7ouJFRd6pgPTSeFSTwmhlnWHNcrvnaf4
5gN6FtPRZvv0as8+c2YRpx0Z06qevztwYgvcd7bZFqOUlV2knYn+sG/BY0sVutDjU1NRRMpQ3lo+
BpXRRIJmkXkqBl7CPls88vsiNTaA4Asz35pwVSl9pF/RCQ750mdq0uGMRLb+NsxV4iDCQ5q3AQbD
tlHdNEESHYdi9aepaseLa63MuN2Udve+3om/6pRKqXeAY8HnsxCcA1ooBI3a10eDhLmWXuUP/CAt
Ydy58reL2OOOP1F+7EUCnFqsCfV8E+XNIjgYEKw+XkO4t+xD/43beiADcLYt5C9OKxw9kEsYqH9w
vu7exsSOXhPgmzwWBWpcFXu3WzQdhVagTDNiVx8UFmz+zQ55+kgqmOv59UjnV42zzqvQ4BO6FfS0
uEL2orTwTiG1DsOuqb4/xD4VIBmKfVWIaNzloMPZAskCxmJHgvVdshGO6bPC8ItM21DQq86aF647
ShAJ4IMpV/GPVuUHT35E4QKdTQmI0vj9El/DvxtBomVhJm4DoM6VyVkuGgUUhL89OqkLL/pKIEtU
we18f6aJ7Z7SERXv/jQLYeAOlhrW5lDPWALaXQczXLMPp8QTb8OS+HSaKyI1EJ1ZXeV2iZDYuFAB
DP+fu/u2cX9kwreKQL4YI8Y+7Z93HxhFQkr3H8f+W0NytPG8D+WVNKBHw8KJVC/MVYo8FM8V24v/
4vd1d38TcVmw4MqeYNL3qhXsRtNusOXTo/jhC8cVPtWHypyozsa7DVJY43RnfmyqKrB+lkbMvJW2
hKcdRaCNPtlZkEk5ddU5tEo9HFNT53ZypazEXRC0mgByNGAZWUbdbsQoXgKHvLFWyDM3le1kPywO
HqtzuGU7Y7gkEh1uT48UnjW9Ov/aVYszQaWEYbOEGSXCKfOR/QXFE+S8DwS/yNOb+yHbsRbRXA5C
1UIOVKxwt5PkC+rdIAcpPiA3Mn/Sc0xilskPmp8ojyQqHh3DpFXdtVS5KJnKpuNyJZGlHWSk+hmX
zrfes0xAxFE6MOJov/4cdg7IGbCbI4Cz3ihVqpk9nZ3nUn4b5KaEL0Ti4dlw+5wF47ZLcrM+DBvg
H6u/kLLp/9gY75zu0k4LM9s7bUO+Nf6vP06xdQy8jm+EFR4dZDXZIaaXkXOAUvaUCZ/wXiqAX6if
TZYgmnE3FMGNaY4eD9LyIwot8IXYwLzf6ho/Qcuu+CfgUMixxHUqv5eCQEJJ4AflOcKJRbQBFoR9
woTHP8u9kyHIuJ8RS8TfGOuZs2uhOxmLmfEaNCYfljGoNKGipY/P1I/K9qEjt5HIlsJmrru6sQtM
ASbgl1KM1JMgVMmlI3l0G84zpzOt3wAMgRdonsiGN/VystvvzE256cLj2A6k3E1bzVeeJrw0CuSW
pmGCqDq9KSdnC7pK5n1qk5TFfJUqbrWlX7qOdD4X+Msf4jK2Q3bnU4D4tk1kM2Sq88J49VqruN/g
XXyn1O6jygVLooFgNPY2KlSYeaNzt21tH3dNI5quGKGhvhvzGnDUZ0sUPAhYvaGfSGuZHa3shQB/
kjxgyeKbsfDrrwmd5NxQZMWXd5PccHtcgBEbxHv1hzKplLOSDeXzeVqi5HTRH5GGjoRlXWl51Nc0
s+KtPgln1X2spkz1rDK2z1+rB3jPrN8IBDKyzH/O6Ewo0WjSvzeHPctXPzSv+HfMJHc/9KymMz70
KCxp+9JmjH0JkBaifGKY6aA/rKpp70XnL+ZYjTizNHaod2Kj5tJbCsQILNt9NKstPtFCVzX/KW11
uFLQ99e5VdH6R+rJ0ofjCq43u7ehb7Wgu9TtVtq1pVuMKeFI1xg8Wjsnq1Pbad4RMPRjtEXe0cJf
aerFBygWe6i782dM5BfDec5dHkAlD/zZWc4lVSg6hgsZiTItiw7fQpRSVjkSeEYBp2j7h9te79xS
PYl4nHFGUP0K3t9nq8+VUAsmmUfgn9FtOdlClewr1tQr63q81YyzX6P8/1MrgvpO3ljDfA8Awk09
E7hZFXnxTUrnDzAAcAB/y/rBzfLMxECuZF9lhOMN2pwdPz/DEViCoqFyrCqHCbOJhiI5QbCWoiNi
Fy9j0qZTRtg14LnoNBlNN6rMHpXk1W2bmIge8ZVgQQq+xKHR5C8EzFXsgfpDHmtgeiAZzcg5Ry79
W8+1jcom0iCb1evzV+urysOa/adlnJ0udpMspA1cSaZ0JURXNpiiLwU3WMWejkul5NmlrusejUKX
USmnbErz2RX71p66D+F9y1KRZTycaX8SrVaHI1Kp6gBWL5Mmy9nfuAhSYYt8uz7lgd4dxQDPEr7x
5YgQglERKVZESy+L/u+Gffz0sB98xI323+6mCrNzUCXRdYdEyBKvBrQMyXbP8ZQwpVZ/mJoRA8CA
LPbktPgTRDy2INU6pk7NNg/O5thzfIj9ggJQD2aCQZyeWZDFfh3g+wFoL64zmdMT6HLRptBSLVFM
8I8gLcmcfd/gMFeFUwQt7Hqvyix+BeGc7WN3+7iBQmyAH9y2fet1FGcNHWyLh+jNxznJS80nVG7v
i7i8LT2msqvq0+nn7DtaYl0iIEdjm/RVY1yY6QNO6jNhJ72Q+uWswV+2mS9gAHyon2eMWXr/V7VJ
RoIhZXZcpT3QaO/m+Kb4cjL9lmHo6VdylMj2jufZYDa3Jo5ktEvkqe/uukSguNuU1m0ov+f//2Uf
AywBf4c3UWWeZWLEpk9zAQOqtMzGMWtoUdevpgcnd4k1bie9hIfSicnGjL5Uob9iHjZiqRLe3MWW
2ThhcCG1lMYhIf9RZtaTkfTQYHI/pFcDmwH5cNvistOXdcPgLt9Yqya3jW0WUbkYVO9hdj95zSnH
CjS0Y1kVyuuqGhuoCHo7aTG9oWMcbnvO88hHRC7Vik35rgh+EEM3dR9igu5U0FyzrM0Jt/BvADni
Blxn0rziitBDVhNOZoFegcIL+hv4TGHsByLQHjZB71vLGy6t3vsDAeTWGB5yVC9GaMrmnT6Jm46h
5GV0+2ssgm1y+6jCOho0IEwZt2XoIyb6Ty4Ap/9XVtVE4DXZs6w4zgoe1a6oOkBpttq1kqLA8Wam
myb1cMSy0OU98akuuCsA5OHoEeSiF4uPxHZYu0CYf90wTuVKNSzwEkaPpRKYRCkfgTd80+ZoV0+o
sii7JB+2lZKfdeHyBXODIIkFRIqyAyGp02qhLAjsargOaiDsMWbPjl9HnSgbsJIZbRtYGcELfgHq
lhRZT2N9rHyVWWVhck/IP5CKi0vPxkuOQYy5jwcN9a6JGjyn+Px+LWsVo79QUNZmSduarIXSEN6Y
FlYHAIPtqWX3QfA8N/4yuTD9eo7pDNGfMM64bc3eMpMltR2kSdVQUp1tHcqIN0cY49VmUtcVaskg
55b3FHxmD9riHR/5YrLd9wFVYo0d92fPmpvgf9Rs7MoV/oXKATvbplaXw0WnbVzNtjtNxkLT4sN2
S93vM58aHiX1ztQRPWj4AX1FEHIZhO31+GsdTp4bEVdCh4IEBWyghj2f3W5mKMjPU3JfJnueaZHV
lNwxiDRgtMXf+I+rA3WkPq+WGtLw5v/5147eLAwGjR2VGDi6PBWRvvfMxr7TGNppxzTbJIsaEX+J
FBc9WszRUVVAnfFya7WAj4Y0wTYYdtJBJAr5RV7s2Bv8RPHeqSg6wtLVYxoTGcziuEubFANPi/XJ
vqNG4DBxv2ZYZMNb82odNqj5flomva8wOs5LU05DNPxj0sBYnqLvlfVEuybIJ8H1dj5PukfaWMt4
04ulqQNh748ZKyFqSlMIAGr7FT3f8b3SdPmrLzFHAGJqyMIxqb5RzzRdGBtMMaiyqvYel5YaeL91
RaswoZSC9+WX9GKyuPlLvBx8pi70hLHi1QG7eosD9XHC97RWsYKavl+rQN64V0kmZjIAxXfFjTO/
LsmWllH8i6IViG5WNY2IVyqgk2vVYSIezvYIj2JgydOaOQ2sYG3QitTP9F9r91h9POJ/uz9exO2z
Wz9GVEK201B1qFDyZcWZRfdJpqYejuxdGc9WtEnvIJBBEzP6+kbIUssb5XKJuz63R7LSxU0J5A8r
EV9Dd2otNTcrSL05NucYMkuzijVWbnYAuwlYP16xX3o/cflDEVreRbHvXGUm4qn1rpdA7tdP4XAW
rtzYrOv6OcU5Y0tH/YrUcOi7ETOHpI4T1kXc4gwkv5Qejgcrqhmhl5j0SA8RjL1WxD22TBu+9VAx
i/C7peCZdqgBEwHz9ticSWi+l6KUxHo9P4TCkjJPt15lwV8968j3Syp38GsvOMTgujLYzYAoKdCp
gokaJWjpVL9KY+qSYxHTbwaxt2S15lQ6JUaet6M6PxI7u/kKchx+lvXIlc9AdNDruAiL/HDjqqCB
37VI5hGlNDcn3KccUyNSUov16yTXD9PRlZNjWhSK6RHYQ17Y591LNQZJobMMLinJg03IawBhD1XW
deG5ihSWtiy1QfLRM96lndASixVDBNjATCbU2B+uvRmFb9dhPPDMuzGiBo76d4y6HIknmVROGvE9
pm2iCEpJej8xIOjsi4kRN90xa6MRZvvhV03Ig7EfyKJQJ/3h0umlKMl7RbYIXcfyJX4OFEk638xM
4FaJIpVQ69RraGFzKWOh9huqm0IIiF6SGSFzYK2m5vJg/qi8MzhpTsCYQgcmL7x+BspERNWgBLBW
0So690JAupb/BqTfVKRfV3KX42E6brLwIZ5IOa+LCqF4+7iIPBZVUmLnodFDDsBXrXUc7/ubuQgF
tODST7e128R8139thFM9sYa/GrBm4hLWLofHbqxjw2M3yGAA+BuM5oiuzNpAU4RLnQ0TT08E1FIh
QJTyCKiHV4XouixBbn1KI5FJSI2VHwLQwe1V8QYcQV4qZXUdVdANucea3Ei5Et9xhYNwwAA5w9JC
K86CbwEiPIP0JwS/r1269rjIm2BZ2RPzpBtV3joTh61ZqoIXIqDX6ucz4FBshOYpVIQAK7+3rB7I
a5dg3TNyVYzLhtz6ONpO9qTl7s8Kn+Y+J01u0ojhvapUjDcx3Z0dMSL6E2Hucnim/WOAd7qvVWL5
ScqWc8Z9DZLQcB3s15BH6uC39igzjRmNg2e3cg6q43WMljVz5cAwjLAF0cZaemBMd7ZSNlgAkD33
vzsHUy60E3jgDYiyvK1p6ert5V9Si62qSjCyoiVXjB+IS4FlCFJEc4AtGKW9Gm51jGAGCbMKfNmA
1ZcP/6f2QH6wrA2+pSB21EmAdBOMohuR9WXX5wj3gJafgZU+6mIu4KTwvM6xP+sft4UtuLRmw7SE
33uLJFeyOnlp5m4AogpSDc3dNfVAQjmqShayVoCgxhnZDXB0XalzRBU/gQIuAr5usmNqGFsQjh20
moZ32p7XWtbNEfAB+mOmglb5BvY8Q0+dgS21bq67emNQ+du73gO44Xkir99DUz3No2k4jkDB9cWb
DZFe4jVPgybqMKDpyzypMRfkxnbl0FGqIt3PigRyfa/0ux2jF6CSDkaTmXmvAvprPvpVDhV3U4Wk
B0b8CiwuqJIcGLAqVQIZZlQxI9kqOxvn3tpE2Rs88NGq5gWxwsH/lT4YJ09GLlWElXs1ZeylZULz
TAUUQonDtS7yPQH1uXdR7PMiuftLittyCmsxEX6CMZJm9CK6BvWx0HQqAdAYawaTVu97ZPgSFKhH
UT3SVXjUswvgg9PhhtykptkdwF5bFlr8zwtvoBGuK6ghaCwIRbob2f6KuOOHTojG0pGSG2ZOPP2s
cg80wWdiSwe4Z1tSS47umdXcYzb7bBOrEOYdgqM1fObBJbaiFkQGiVNEKG5qo+jO67k5/1cVNuCK
SjqYM5HV56Kgol0GR76LYtKx4czG71GRI1yZszeda05v98r7Hkn6SJUQomsBIUypvU4CASaWQO83
Nz5RASz5gbfXzxzuRjBuhIAtOnyOTuU3XY9UlEVbSjRtV6III6E+vXX2Ue+iNEG7FHNFl49JItau
rBubL6ySSeFVbBb8r8rj1okHdePncH+rhvUHcB+3QebaPPz2y8m5eZtjzDC2tBntmmIPQBeyR6pj
Vc+pLjANzmqDsVIccQBwpZBoanP2AaqLAkZFQaieKcNcBD1uygHqlqA75lPtcCAk4tO228wQfium
c075hpaGB3mHqSir11c8xj0XHR0Md38iGLh51l33Fel7nKmLLfcL2jErPwp9Ae1wdoN5jSPqI/ma
ZZnLPNq8nv8laCg9LeQYEOh6fiCxPAHPJnFNP0YARM9cP6rJoKS8JlaN0eq/yCNYyLY/oPfTvgFZ
DdNhcGb22mFJbdICUHlnARectWMhP385GOV2l1ihMkqFhc/9ZN38Snlpwa7lWS9QpdokibwDLTwk
eU7tAocUzXiJ8IOGFwsvoQEMjcgqpDuTGVEBdL4Q2a8msznf+VrIF5BX4Wi0ORLgtlqNr+j4mrS9
oDYYz8U7R1pO3oUaQYk/e8R6Sqr+AwHmirA23QNc/PioG3gOs4mzWtwPGFTLiS1t5zH3qsL/tq1o
pWMbyW8pibRPQEKP64yLOmMdBwno0AtUdsXhyyKBiZNcThEIgKO6e2QAGpy9Cl2ioXNVdhz/hgWv
EtF2Yx7X+EoVkmXSJO96Zq8B7lvrrAqEJncY5sth1DhyrNoFBm3zAMMDVYZC77gT5yfPhrdbxG0W
RhpQIIMKXLBwGZbYzmhy+e/OZfJlDi9ApaHNC85jiPjuaG1wODGoEiE8+B2nEFSLpMmPub9N7J1o
gTlqynRt7eTJNn63sE1pr0z2AFAaX8MQ8WSPF0BWC2FHADiT35GdoqPPgm59Pljtj5eXvb0p89Xn
/x6HUEcwrEHb2MwpbG/TDb7XBHXAgTgQ2ewNf4STXJXYzeyhi/AzcdbOxDpRWAAMyLjOqRNJhEHx
TJAPKfoIT1xYlRD/3knWpLvJjPFnoUR7w1SBiF96pn9PLZiC+iFasohlrjUA09QvdFoLK6tQZjdL
uRXWKJwqAcFeP6umD6I5nFTIvKUoCBKcrGHb5s7kxPQA7QWvSyrXxtGz6ajP9doEjcTGk/tEsdEB
DDOthUeFC+3Smx45bp45AWlTTXkESJRQpbtsu3BNJQhqz34WQgFZG4vJXI3t9zboO6bm0auwxnif
SDc5OcC2ZmGzePUgRtxKDnNDnOD6mrayv7Io3fKeqffGg/OlBCWrE6uPHEbiuG/hYqACyhP9jC17
jI1K8Hcn9/tab/VxQO1KLVvmBKFmobY3KzG97puypP0puvqTn+lmxbIelMWMU3TP9jzPpK2F0Xdc
Rz8+uz9ieXbwGqAuvF0orNn/bAo5JCmW+WfMNn4HxHn500aioKFbH+HaF+t6RI53cnzeqS4QL6o8
M0COFjfiQmASwBpbWLikwuBo6cJ0N/+q33kz2dmkGdIh5QNmSeyg4FPJBx0dIb6yMbmT19SkDcNb
/OnGOOWUX60TwvI7M9qtlV+sMU2xnQZ2lL0xFtoocNP9mrY2MBOQS2iSXKBQTrucdkuAL7YTfJqY
1B26nA4PrAIm+xSFeAlhyxjz6irRaF1tRk0997EVn3+4olnTR+uabJStu5IeA7pAAfWZy0/Qmkrf
hApptG2cGpoxWZ7di2J6VXtyj97n/D+elbM0XL6GMRSxjGy3sSNddQzuOYmNgydrgAz69Umlcj9L
6nF81TdtiKHL8e47zlSnaxxiv66XzizTy5tdsaEXYvu9YY7hql0XG7+QCMVjfv02T/esRTuAdaGZ
0XpzLheu7KAvzawcivCnNxMTBvpth11xCUrcRaF99wFyiiltubgkvaCCtZA2+NhaVfAV8ruRoCSL
1KDI00MkgSzx4drHx3mB5BohBcvZ0J8uEN03lhT+mfK7gHwaxYAzAFehtlz13SX4g1JAAyE4RV/N
jd0R9HTi+xmm6vsPxVO8//LfdBtswz+VDupcs6ZZdCHyVZToDsIS3S92mDPXy9hez2i7ZaTv8JtE
RZCtmIN+nfmSWJ+c1cbULrC/tRmmo5LMYnL6Q2e27NQKoFq3ERUxSNcYXyiwcx9h1uBP2httYwLc
hsqXEnWa3YQSNaKr9yLGO0BWP2lsPEHGrGB9B6y2PcbXTQ9TM2Jqre/SsfZbFxsq5SqkZTzRjFiM
CgS4fH8os90AD6VO5LUx0U5iW7Gcdv137lPIVQ4pIBQ1tUPa1IKn7aM5+slpN7NUXOkw6QrUKVHm
bijz7Nfucd+D2p4OrOWXOACg+9Zpq9f94MjBlCCcZb67P6Av6fWrcprH8KsSFsc/qRl9P/sMgLTs
m1MVRav9PYo6MZ0YPTKovHWDwlhTMdVXwh9iWQj+TG8l1IE3pHQb5yjR+H8wWlM1sRL3gniW7x8p
QYuesGMOQ6ZV+1ECglpk8qP5Ge5vvkOGR/ad4gnoeyLlbCU7yj1IfvIsRxIEALT1yT8eyJkkte1S
9dBpT7B4ujrLHaNpJTDSg4WTnMIUM/c3x9OR4IYsYamHO4Ju1mtzsVYMOLgee/SN7ozXBcYMM7CJ
ddRUjp3jst174/7j6dEE1fYP5K3drtepOpuGXGA57/Lm30WhQ9Pc8eFXSql6JXUtXfiB4eTBwWLx
riyxKMDcjDHIGfyhjwXxFXlqlTHtiJe9wogRKy71qWeJQs5IZ5U2YYMA2UchxDoY6j0NL6Zi0G4X
H8wj8NDidCghfHaw3zjsTeLVaGwBxHSOteNstDtN9ZXsyEPjparmdoxKsiuEuG5JufivvvvvGiuf
RZGuaAN5X+xKx5BvzmTBrlTICdqHNrvB86qM/jOSgh8lmSyvx+wXkKHVEfYZ70rr9OnkS2Y7axOr
p+QIJoprl3HA589hG0PJrLRhpsiT7o3+hj2HSoB2s4DqS6ukLaQdLuH2uqEgQRJsdWvxZVv2dlUN
ThpRKM1+kW2QSmCmHCSGV9yqV6HCxZuNfFqiJqsiXk+wHqRyqOW6fE4VRX90cS2zIF1kPQhieGjk
NHdfmifVfdTQNljtEvhC6KGwTASr2FAQojdbO0yGIs+E5j7p4PfX25MnkxDTzIDUb2yxf5FYobDQ
p0XwznBaPCKdKN5gSM2tUs2xG8FnStzNw8ehbaze4f8Jyjcb9quMkk7eOoMFr5APRpgZnhKvcIkp
hlmanBQFfJrjZ3DtKzx9IDH8yv7uGbDzvXQ1AZmv88KYEpuuu4DuJbTJfzMKHKV+YJ0kOJ1TAucg
BkhFMuFsQt+Mgi8tEBJsk5WNuqQ3KHgFOadWyAR9wHsMKXoQZODb3Jva1cyoSxQVdpKRQEbFpUOO
PWetEoG1BZm2JV/khrrDIwD8/RBfSBZx0R+xNOzuX7ffTqvEgNLLnaIrmHjOEVHJrIdq/7+QIgOZ
wUlAfMuUmsKQnXD7VhqeqdJj8Q+2pjWfpAsx91iPb7fC4c7CGzuaWsrJZTCeb2fQgzbItCFN6E+p
ZzcQH4UnWoG1DfiTDkhorDzfQmDgCP79gCY2BE8Em/ce5FZc1kcXETi3OFDnE99wusUGtZjgFRfa
aYZ8BcYWxbfbVe3uVp8t74DcnTZOwm7iaj9ZB5NGHZsktxWBsUqe91rgvI606HdHHiFVhuVguuNy
6m7b+cSBGkGlbH7cXsfLnbmMiiLhZbA6mRX8npZJLR87DBcAzKcbzKUQPgb51Y4bl4MIKnLFTg5u
iMNT4CIy/SJtnG0J/MpjA39cXhuAAwXbSQ1KLnF2BxgHUzxjuqWs4CUaZqFXpK7gqWI03vMdSspk
FE0OQuJoGQpfl7l61PN+r2duB2efjgcy+aOH48NI+cAYkPtm9BFwDQ+7tdjiMVP3JvF5nC151q2c
Ge8KfbJNUHxRW6Lqs4nIqcCqoKligZ/c/lMrCiwoU9edS1gNd6k/ZSp2FXqgzqR2CX0+Pu2rijFs
d+AqNAc0RUL5pqpFVO6C7C7N8+04nhIEoB8h9TYeYud9mDKSJFeheWCuucwPNYsFjp5tc7irTG7D
gnl/SPec6dkicswKcaOUBT07pnr1melXd1E+8gcWMpNoLGsawwg3AwYNc1CDfbEsjFNhTbfsQDLB
gzteWez0ELBqQTnCFbuXA25ho95+vKe/DPYB/TlMXuJ+KjqKUZXV2OKUDJ0ajMVv+3uoFHmKnaM7
VSgbhmouTVa4F09qiEao+bXJLnADCluoWCBN6vgVcO1J+MdbWIuPFfIip/4XanpzfLm8A3rXK7x7
t1RHeZb1kz9B1fMN8q0K36gaBVgDZW3Hs+BcF4n0hm2ROKNSLy3lMEiBdXC72usa44n+met4XtEp
tTHS9ayPzOefDqjNKFLIkntaEVb4vhh2I50FvOgk1VzLuiXHWopsLkxykATKxo/PqqvBFkZUJDmk
wzX+fjJlXAWMKt7vdj22/ZUNKKnBouCwLNNmuD8EuBebNM05geQ9VSpY3pu5+9KP3YaBTB80PzYv
KMwBFlqxBRF3v2Xu6dqPP9jDLYha6vZflykDl7F75Drt7NtAEnV65lG3GkxX0nBjJSdznvlcCux+
YqBSlGhZzRifKN1KqmPtBnykFofvrSIcOQFYmzwXhcSCWCROwsD857ELb1olJcTiiXk56p9a6JjT
3u2lGgER/q7j8I14h52q7nMvv1z8uJdW9U0Yz1qC+GEYMlni8sGZMBJpxxfk2G8NG/8mnxTwNG0f
RRh/7ES71o0q/mhnQxvOmvpDzXigQjxstRbUQIn1NZ86e1rStj9ewmuEDkQ5b+ekYVwShig377Ip
x254MxUD470cgbQp1qJk01lMb9kQEReJoV2Sk7GxqJtwMxaLiIOHqCXvwJ7wAP0XCyez0w9ShjJR
LijIBPU+lbWgdZxuTjzZ07/bKJPDzxNqSY4BRZQRTm0YlfO3ROAhpu7nXlhWnYl4a85xEez982Op
LECoHXct2wlmfBZGBERlyOKsKignQ1QkJ3Fn0yFwOT6sEczHhcbVx9Ta1vtV4UFYz4sksOHpBiMV
KowqlrDg8qIVwYhjjK+qM2yG6Eq+cmeQ4UsCO3W0k11YDZ4lZ+4VfQihcf4X5NIUE08YsYpJj2yA
20gk7tQ4IHVSp6nYbess8yCrbGO63TMh+xQ0FsWB0nk3wc1G1cj/gorrGLOtiAwAKcNo8RwitH4i
2FdouLvXSUoRwaKLoIzVbqJnv5AvQjN6uSXff52ErYpRrKhVbocrPWc/tIImeP4vK3QiVX6GOcxx
W8LAO1DEkAzGvgUIE4Z3PjiqzKP06z4zqz++tKsITAHC5SlpbWpAmRVzx9EvAJPQINNU8D+zUYHz
Yk8TaEshDIedbtFmzy2iqD/E4g8M5ATMn7fY3FyxiPngZLwxE8GbS3FkV6J58yGtPzjnVLRxgRdw
+uSusMCYtgN2wxf8wEHWkqrcM8k4mD5AEMMp7fpt3GyowRdpGpPQJiH0MeGUdfYZ7QAMJ6vG+rva
ZeMqaxRmLMFhf0FeHDA/fduTOxiTwKXtXjC9J9fT+cSI72S7RM1hAHroUQMG0hdvvpGwIrtpwZQs
iq/gJZI1BuavWQ/dtl+DsvsMXezdN8fm7KH9PJGMxqKHrbYEkIl8MYIcto2IORzd8MQfVQCcpM7L
vK2JmujZkm2Clc83r83FZp5Emaw92TMpvSoPCho7NAtmjmN/XtG9seZNUg8xCH1IU8kvNT35JzGz
cO4T1nfeRzkhDToF4xbHRkeKjTTfGA8M4f/iexnc5NCnzJdLM5Ems4As0ZAjDqximWwybZwlB7VS
gZJwxG0Dg3Q++o5tkfSPOjSplVtLU8vcF/VH+B2yt3/9YDAuzdTTmZwh/Ac9v5r/JE291XeURhwP
gFI2Buv5Utwgh091rSd4AH5Fr9BTNWpSFg8nynre8ojIJfPewy+4cC6YAjdEh3pQrFiVQ6OoKIyo
OcEEWvXyYR3RaLsDEbElzNbOFaDMZgw42uqWK8FdsUBV5MLDNwyk1DoXkYfMXaRDNxw8JXvhNl+S
22jrf1E2eM6wY7god1LSx6yqgKGhWpxwrzs9GOjmwGOhZc9WKZt00l5qRvtjvN95QoLj04bJJqcJ
3VXdcrfhTtytZSNcAu7LSYsel2trMCvJh1dH7e5Gi2ZYXCm6+3ad2S6Kwuq10wR3MZpM+bbIZ1Ww
bAIsMbsU7QLBGmdQlvWoE0c1YhkyQvY+QbJr5d/Tjmv9MjOOm/xd2inJVMenGbpAkyo0ziYnZRF4
vUvBIlOXcTtxWYvoOYcpQtxF2HxWwLh2uNnZz88o7WMQnd1yzJwv/MQT+FhJWh/jXSzX+N0fVRzc
TboNoQgfNRWcVYzQAlzhMhMl6kw0sHFGODi199dSS2xJ3ori8LiSfGy9TsaBReeKYk3egIqz4sh8
6X0VcjSln/0VNsYHSRutk5pHvRCxLnnmPq4H+c5UtV8d9eKspiwrbr/YW0zzL/UU0jYcwmDrBxIZ
TMPXVjyS77+ww++yS0FsaDG5QVtxYJMlRjWXBUDZavf/nfoNAORNlGva57xT7ZOsv2K920l9pqpy
2pxBCK4YMbLpiKYnRMtMhHQytUHnZoNd0xyYhIn2DGu262Rl2TD04gzrciyNYaXZh2+C2/49Yihn
SiwoZrYpzFngilQs30xzqjZwSI788o92fpBj2L3JlrgM/urHh2FrpIAtytEZAtCRyk0v/enMavJ3
cyOPvqGYIjIQ8/Dxv5DEC2Oce3TgKOln96V0uU3MpO0VJ88umc3AMP7j4IunkltPl96KdMjW8GMX
RZ+sFaxsgtUACzGtiyTsjpGBMB66GnS37G5X1lo5+J1P6czx2Yj8SyNRp4DjvxGLScAufMtxmuwt
fOPvNFfEjJ2AIjScj1jGXvX5lTEe5L1KtuYhKsF2HzempfX3IoIWMSZYTXfN8Pd0HzDyLZTVPKPH
v/KtucxG/6WIiYLKxdMZNfudDrW/fDuh/PInCcnINC0w/R4bIotk/MVRguzwp+y3+AToze8Sd+TU
qv6tt1xgBzQxBG4eY4df103s/U2+ewo1IrBSzbT4mQcypjKjuojizc8cyaPKPgVDoIE8s7Z1/6iP
CePQNqikFHuQn+ojyEqmHQ/6sihCsiily35kinNNzn/dK/xPPzpM4wXWsDaWOCIHCacjw3V9f5ij
0G/bWokOS2af5oa7c6r6ldSgNHokB6gMFL8u0UUgr5JWje+hGCirpsyWbcQfBJrXU1+Me8TR4UWu
mWUqm8ahi5yMpAYly9ajeLlJy5MzZh76LO2l9q2Xydx+J+vnzMRdhI3qQcE+PJXAAKK40eJoaFR+
5oITQaRz+Aryyh8Pw68167MIsxdzBm1jj04vhwWBmFT+YvQumabmyl7FQgPT+Q0tRQnrhxZYB5Et
FeT4T+vDubzDnNPYmefsl6s6BfJo2xcEIRpITCPrXLzBxCdv4TpQicczT9XqMNHdUKCunTv7/2Fp
lhTogj9Mbm2C8n/jxcGuUe/UE1y+DFq8Vi57iuRcbTdarq8VJvPfFFl9P4nl1niOhJWDLWUz/lFl
Bb5utOqZsN5um+ORo+bm3N7cdIzF5Du6gh3TwV3aO1rZx07I4PtXYR86Ti/oSR7g5D9ZrA03Vpx5
b8eGCsuB8uBEeMjUuTI2l/ibB9Em6dqChkSSsA6lQLJk7WSBMf/Xdpw/Bx4sNqF52JnVcFAlVSxx
bEEaBSvnzxGw1xVaSVxvM/dE3J0g9B/SDXVdmA/OLGbc67mRTkA26vC4J7ByxyDIBv3KjbE6xdua
6N5WULx3GXpnTtoFFhlvA3p+9F+jcYz0TDr2h1az3ZzPMCkKvBkyeLfBq7ErEMtLryjaydE5XNY6
uzAuheJurIAjNMCut2x3LDnHEincMcNk++SE6Wrmlh2oBfvqngES3uVwEDcyPH3sgqKv1apVOZdG
NrmeM6xHKGVyBIsWB2FhsSKzzM3FUMZuUVeV3LvfH4qo6SY/QvC8dQC5ZlHOXobdnqACpJhURp9L
kdLP6GMOYcMblIk6AERNi+iXh/Y6b6zSwPeoFG9HplozHNbRjjf0t3WG1ts3l+AxOlZQVvpsd/2p
Yrynfs56LMs0hCxe3aTfXKxKY3y316UjCdlYOEFul5jaAPrhFYBpLNbwNO+rKqsCgW9l6RxJbCiR
VpPED7ANXZfdqePDLOlIDsBqoZ+/LfcnIhELuCcq7vC+MUErkBl0zyMxCJJaf+1oYv6O80hR0r8d
7E4h1SblonViFqIkEqYlzXDKxN7q8ywMVuSKoVCAssCcz8f/LCS/SOYt0eHSemAfCvBWZn4BB4NP
/B41qrlqdHd4B6453A4I39FF+4yxCf0doxs9BAg+1OKXix8XPpGsEky6uyTLas7CYGIMtTi4QbAV
FCOqKBV66i7/a2wjw6iy8Ocm9j3tmNVnQwXJPJZYCu9cbRLh9de4dkbRw5Xv/BTID9vnfgOUVLIe
9E179CDFSb9mWrSzlRbkp+g8kWt1+FecUuqfEdbkPaU/XWVu4Enn4UrxfegzT7DHDwMsBcPkMPCe
M11fw9VtyST/jr/2RoMndC3JFvrkc3AzomMQGjA3iwHdDeepV89qduRz2wWabzn35yv/gK1Meq15
+/i6xwa2XwIupZxHpe/2vAHYZzLMgUB+hBo6R2F+2zK7YxiDYaWz17BOhkhGkbW7D4xFRA+Pfvbu
IK84pa+HoyNFvm7D35IP5DyxyXg8HCBtvWw/qsFSBxaj2jp+1qvET3NnHqsbMGExc2ybcucp8uGl
EeB70n4jF4mhVk6nR502nm3qqdUZ2rjEQG72wzfiLUwNNrx41+WlcCflMbTyYIZDIdOcfjiqGCz9
Z34oyLXFY54OHhBx2JaCCb5EbTd3UJzyWGTIJjdet3JEIH0uCopA7r3ejgUhj2sxmmL6YRnV6/ke
pHH0TOsuu4NToLRpIMFkMFzYoNJuLfXyj6Hw42Stvt6dx+f8uB/5eFjEwUQhea+rhBzQxs/5LaeU
aowplWJXacHYgzkSCsGl0YwMrJfX0R9gmNylkBEKy7G33wzDDIyPZtWoN5JX8R/Pc0f2waCzh/8W
7JCyvxyfeLIsrm3nqOyCh2K40qMmzRvtisNm+RwwxwAyejW31uadPpy5+zQi6ON0vW/hLcmVBrTt
CnGDwez/zEWTqdZoRewcW1keSNwzVoZ2HoWA6e5bgcPIR67U0DzT6FIHk3w+203P2yUXm+vWDyKf
5ujk2Q0szQBAdBjxDMQTNIfpwwjewF2adtcPQ1BZZA/JwepPVPxIca5fz0R8f7Sa6U3SWSYqY9Ua
tK+uKgpV4ofTZorvGYZom+Xno+sn0aCBjP6ZfeqI/bkcfZQdln4hjnJeEtnU7JSn83RjdXPtVfA2
SFHGflBeWEvR0merQpe2JYEU/02Xg5KkORkBVqPYyxA4n22qmTUDCD7Sy61PjMO23W3vUhcCC3OU
xmLHt74MfY5DJXOp3UQII7HS+7a6ZQRUmlnd/cDGNQZQ3iNam08oGRZsnCIirLTko7UpDQFPc+wr
IFyAawtYCJC0Gc/fb6fCCD/m+bMcCZ08fDq2VdlYkfDdv+4gcpdXJlcsXBaGgeWulRxO4KpDTsfd
pTh+kkDKEiUBAtuOAr9ObViyg+gNfJTIv4ZUJ7vJAfGJndzWLxOlK8CITANHDUiz1KzzGLXprzK1
UP9WN261ie4iLZopKptF/VM9+RZs5kMi7RYh1wLyL1AgiymcZPPh4EPqkbja28kw2C+fOSIwjt2C
i7B7N1F/PO80f2PBh7WST++zeq7JXB1QqF+DMm4tFFC9kJgDSNoCJ8FYn+wpEZcVrzsk5oltBw4Q
m4pkfh+zGQgEYWgNRhWEfjGLVn18PrcIucNvlOFVIMc3a4MwlDaT2u+fSmCkrucxb3pK6QwowQgJ
pI78JJMpdvMCw7+mHIFPywcldKuGTjHXorEggmDNWlbTvp50P4/yxIIEhhVX9yVAs5OQz9QzxdhF
4augUHuLc1HlR6M5rEC4Ofo9hKB0vD1CPTqPyLqNX71FpiMYLEMJ+U17U3HDJLSUxQBi+s6l+4Dv
0hPucsR7ZNJ4pyZSVQ0RKORCNYHsY16aP01NTQdKa5YwiqzPtkXXV1tUGakww7iTrh+XEk2ywTey
MN3RvS9o7FHrN4JUFCXKS9NCYOb1U7F6Zd/6XiqrnQhPVaz9PIxqwcm75clYr9lur5ZyxCvdrx/u
B4sa1i0WJdDBBSJNyJZFkaliEHlJtYPdj/w9dMwlwjPvfHcDwO0Ng73tU3E9l6+O/VYWB3gW+zKW
cUXG4GUIBI86injMdl9fI9IT9pLS1G0YideM0Xx890VICAYjYYT3FlmjvqOZ+2EeqOtGyBsXgUiA
Ps7KNXsHhPu7TREKZBmrjeVjGQ/mm5j/FrRGFmD9vqO/vRnwUweCpaoY5SFBTOMVLed0+Rc9irZo
kGuUiSGNxSU8H4Xj1x2vHY9CF2CsSpbXghkdpwWJ10dPWgYvp7vz/cImcR8/eHMUGUD0l+IrtDAE
a0M9GsV4CgnWVK/hBkxiMu5T+0N12AqW4e0J2raKUP1Zj1FU1FWVmihseC11rDRuDFMOt8pqkmGS
0l6Is33SSp+iEXlLq04hcSCDtYkOng3GJSaPcu8DL3pB31qEt99Nmp39zNySUsv+UcBYzGB8HKqf
fvB5muoWa5F+c+H66X1j23aAvlB72hhvuHDYTL4TJjODHLEOJZIUtvNWM+L6oV9lTKudaURApUvl
fZkvqXyEjrsqv55PoFEzVs7/eN+9o8ptH+gZOBT2lHjk6qRtSG+3Hoc5P/OE3k9nVcPVjR9miFp5
JLJcWMN3qgPPP3wezXEWQPlFY9sOBSwzZzhDK2Gs5kGVzjvQClJ/9AGts3kBsL8bwYBfMBKWSewF
W792Zr8gTTnG5Ac0UyuVsKGIOdpa+RdB22tS4j701X8xekq+LLIlhpnScViNELwodsDbTjRy2WWT
hZNMj7ZcgFlMpvSDiejiawbvRDAMhwFC1eGjmkIauMXwf6AWEztHqSItWnUnq/zsRAGSNJltSxyT
NJ7vmAQXygs8FKTAsBrvpmdaj00tPxEcZtGDAD5wbrUKzkEB7KVGt6iyhvIXfcsx1MUNuv5t3GlU
PmxONIcNQoIEX9cdtJrZZzhItp7JvbyPdNx5+Hsc26TPLWLYrpzXceAQMMl2rPMbhWOo8jCK0+BV
PlzAcl5WKTxdsRuJBMtObS8vS085X+N8PBsx/KUzS/8ODNtNnuGrMG6/YA1K4CxCzm91ucD172KW
1tUbayUQ8n4mO7ngGHTYkSg/j9rGYd8ragAbMPPwiKk/uYPIYptyKrN9Jixk3zdX1hFG5ElB3cFx
CR3qW+AMub2FG3uWLpp9zoU4jwdSVNogaPXaWjLpn7zuNI7qVSYU0O91lndF7lMy7/NoVUz7LpEx
R/i0todn3UdM9iMIKtmPmR/v9Qzz5I5uWkzD2AJQcSQzESbFMJsLH9quW/TIeQQJIDkGwxJE6QyY
P/JEhPJp4zzD3p9+H9Y028UeokXQFMT9qVVhu91piGYdw1IFp2rpyS8RtD6GBpN56drUg1rIhao7
VbNKo9Fxa+hhyNqKWKvfEslcTQJto93bWwajnw+YHrhvxuJcBVsW6OLPYTMoFoKZ2xpJHL5t6YiX
hilcT+DCkaJcSl6mEC/M5eWZQvwcYolnRaXh2aJ6BUPPm7K90E3uzvjir/zDE3dsI2JskGehGPi1
UPagDJs5uMYQ3gmF8LXu90001UnnsPLgX2AEcUevCjhfd3J1phLUIDx+0fy75bw8E5T45PYJN3MD
Afw37/nj5L25v2TgKc4ZJYJeIyG0mhsVb0pXnmL0iYAMPLlrP5ckWKLzIRJZdE4NGxvbqafwIRTP
UIMt2qmsghs5sbLCfG7tc6vEM4k/fqnpQeaow6kol9M8dqQ1Cq3Ns8pEdydRzVCvbth+BXg0jKkG
NSOIjvnm3w3gBUNHYTN/jmsscppUwUGTJPxHWKIopjeS2h0Lc52alTd9OCd36q3HiHTTvmEZH2oE
j3lWv7/vZScx8xvr7f51fP1IKfEMaCBEVT+lIQMklMQUQ/H6XkSelZdJfkWssnADkjhDn4M1I+UN
CVDZHlcvsRGGTU8WcFPAojkAmXvFVtY8/6fiVCQ6UvFDHUwjUWQySNArQwD6RpbqINZSahL+3GSZ
KW0Sk+xPQGDXilFrnT7IKw0h7xKEXx/r7mUTgTbEN8GQnoiTqYqLyWvpbvpxF4NcxY62JPUm0v5l
B5aynwHmXhdBLd8aJr6AB3tCyFn4pZG/yOoxAVWxDdubwHYWdf6DaBxfBKVh+816Epm05ZckOB7P
aYNQSvaWE4O3FVU4A7VmzSyxodIcohIcfvs4KYP46kP32f5N36ujk6Z/wO6WKWAppL3dkj4p/9mk
mVpX8U8dY++ZZkszSoIlme5TZIB1qjIVfgN3k5oBZnRhJi3v6b1HtrEmNafOu/n5zu+ySfb+FKQo
xoek0FSWL01/Pg+BGedBWeuBlUUCoiBvcFBmI9RU89M9o/H0n/1pTgvRKJRbweAwI4BC/gKNJtes
aQVpHy2m/v1Y60988aLikGV+G0cHfLktVRzqJG0I5PF3IwNfHU/mtOzwAcpnE7T1S3rAMnpO7FCc
Evd6obK8I+ndRROTeQ+yReZj8TILcrhLrm5Nf+9X3SW3stV6sjWchxInx9ASmqRD1hWRvr0UbVMC
BSTmynp4br/UQhQbw+uTQLGuw87zHnyKUN26RzQNw4qdgPUz0kjqIShm9nB45+amlKhnbo8wKxbY
ltpCzUn0to+NiGT/vVxnPrp8DXExtGqXntup6/dgL4UDXLJddnkJZpOv3XM/eZDJZeKqA092qM8A
Lq0/mfFYkkemnRBdV/ezLg3QKyrhFQL90h7gKYA0Uwne6hz1++fyYsbDefKPndX0R9Ka7Gh9P1Vu
/Fyye61miMgsRtoB+/jcNwbk7gmS/gB/vjDDGf48SnX4mroSUHDVAdxdxnLHFnsw8a7a1+xAkJjo
ly/PigHWyz18F9WFMi9P5NRoJh403zSNAA7TO0p+MQctrbkCaD79ou16Vt6ZxIoKyThxP9P+8pjl
eAWjJsX/1Nl8FSBmF3BEtUFa7jIb2SvERcLWHWxdMVWKG/1pQOjdLYj9kmWuNvjQuaAFPr2Eda4g
G1AD6XTlx3JcIOMQPzHYBp3TyFYBbY5MUxX6QNeN9NVYtiOpU2CT7k7IaBKKjUGrPvrwKv6r9ktR
vHR8EaQhqSFeyPwmt/vkZhj9aJAVAPwgd5ycv+nxtTXmz6zx9SBIaTM9ewaKgYMzzVgHiB9zLE1f
r7Y6aKrlkUp04LwaumbE6JJH/vH5zlguY3C/kDH8QpcS5RfoUXotvn+B/ZLvSAYQx43/fd4y+EmW
UvU6RDIVOEnJXK95eZVQvScmC2s58lulfcRjoxH9gydAFqHcZRkReXzUTLStwNdqaqstvaFd7aJh
XjurWoSi/VGXkXCQJt9ZeFNh6zE3R7TLftbEwIdi+Mh/c55+CpcGo+1q6P8VRQNosv+bCJY/8u54
6iQj2SXNjSPhSCsvJJbljN7JM/VEZs4jp5m13WseuGDgz4ywrtmVS423iKLdJQvmWfS4rlRJey9i
O74bTL6pkTtPvGG7/fQ2L/a/KtirwgZyyo6cN56wuxmwtWK1G+0KhRaYjRmJVFhvrPLKbkK04FSE
3aniAvHM3zzhd6EFVGrVAiCt29f/iBsH7fKoaOtlhHLYsBEOwVzOzKwFzkWmztAZ9Kp2DhUU3Zmc
QLUCMSd7iLwXSCxOcWxf8/uuNP1Bytd7WmhRxKGaK3uKfYORsewdm35BRcCCvfOt4mUoP+rXJ1zp
D55VCNKTDd3BCOjFQVX4GWUF1k/LZsuxKcHmZV4+5bsY2wQj7Ww+QuhfI5BdCaIoFJhqZV/dR+Nz
zJAZ7HDB5djQ6FreSbSrHFgSHvpcebeRyHNP/I2usJycefWtCDDzfJ8ZhQpkUZuQVKIHjJeJ1U9x
Mc5YM2eJ1RSd/oQw+JHn7H+dRngiRihHK5eL9uWuMf16Ivufzdw5qam7L3NtM3UvKYH13wpXxMQL
acVpNRSsLYBIZ719ufFpNOCrX0mVWh23d+09WHfc5b8tt5lQy1DoHSiddIYhj+NUCQfg6Oi2gynm
Vsql8sMRzRe56GbtPpcDY1CQHrbVZ/voU/NtErshh54SB8Zjvc+wzXMqI/DDX5pJ1hJYGvy3WXTl
2eZ8cIAdNZpY//OB2LQ4ya+t5jvbeabmODKOItLxJrpum1iB6SybozGzk6l+UP/8/vWK7/jhXv/C
xss5cYTnXn8r4BYMgKYMNxnffi4WaFn9pcq+I0RCxNCF7sI4LKWvR5UFGxCbAjDz9II9oOgtpnAu
A2KUlBTk59siyuTSeOXm/H0YKyGO8395Yplj+JKVVQvkdd1xCwgds7LskjXDCB3fAeQbaPxEZjP7
tsaXwE8Wk0ayRMU2K23oetJcKfbAxYRh80tOjxY4J5fUK0lo7R367Ooep6OJgMs/ZnTb1am9DeWC
PHYYfja5ji3ZSUX7x4uCkLGKjkEFsQo+cmH4zknQhlxgCI79xpGMZII6akEjLJfuhFlwIhp1iyeO
p0/Q2u9JDjZCHMNkPtNKDZCfGnLum95bGunNx+0wVOKC0GQ2sQg80dD7Q/1Mw3aC5jiJnqRGnIju
cAvo/wgq2U1dBiMvNzk8UC+OTu3DcckP0KQT0eS8yoby/yhbdZDNGaxBOb158bNlrI+qPd5kcww4
QfyDs35OeLZjqCTw88xzIpvBMPu+7uFfHXWSxwPxu/FT5iN65381FZVzDKoUbAHPzTYHXXe/2tf7
TMeSjVxSsUY1nYPHk4xaln2FuxovF/sqT1q/hEztJOC3Udtb4VcB0qV8HtB7a9NDgNVd6o6M3pWC
Y1If2l51B6c1gJm/rgz3N1AKuPmpUoUvNk7l6LxGqVX880+aQTbVxGuzx68Thz3k2EBlfthpLA9X
tuaCYer/wyGNmbUOiODZHyN1gUyE34Vm6evoNpALlslEy3ykVoa/rOJoK81muhz17/tSiaYGFqJO
8zqATsF+gO/O6EeKsBcyaXXAyVRwb68/TBcK4cU4UYSP3TSfKcV9C5ilJ+cLHnIL/NoO5YivCWMy
sQIKIAtpfJDm+sPg/MDSdu9SjPu0rcdJ/hR1nN4jElYdA19vuqmSQRWF/4Qug7lUWU8w5JIs6aj7
0FFRlRgM/+Oo0BFtPU2qnZzwnw1swmu5koUi9IdOU0/jubPzjG9jNF+5UBNK1PwZ1QQc+b7hfDH2
Uby9sSyJgvKyNzFHsmpckKMd9yrM7Srjg6cORb/Vybih9QxQ83E0CfNfG1SWEhIxRhPmgvuYM2Aj
SrdSEtbBWDU08Vk0+i9ElP6k96fadIrrI4pdVZA1suC2B7nAD8MHqFlg8FB+S12+jrL3IYTIs8A2
PcTXAW2PT53a+kJYfLTyzZueF/0tRM8DNLT85LCVjhzYRu3QbrXciUq+O5DseR/8VFIPdVRHoAmx
JIy1UNIphg2hD5eDOENVoegvWaD5aWULdUNBJBnQAoo4OFVJbTGwlc7IsOVt3J8fi7cybFAiRR4H
wfslRnuWXV2Y1pw4jNv5lizEVHPvofPOnDc7a0X9EacigoM8YvFiekvArMFS2cgibsavo+ya873B
DWdDuQzlVozzLhJUOYjZrmeHo6C+JGlNAcuI5ddaO7KqnUhcezr2lQORhIYX16G/uEcElY/Iz5E5
cmXLb91e22dFvZ+Vjd+dAeXYDEBwNcJZ9eVWodKr1xfRe47roV5n5jMYQrajZyG9bZCpRMrTRC83
y9FO1fOh61lZoEfF/pfKfe5G2tFIxdom0+wfZJLFdGhtfGQDsUDsD2L+zDBcNvGiKTJtYLNBVURd
MNC3mWkAOa5BldFcdJnEH7s/VLWzPSi5FxAU6RsViu9rwy2+w0uCMf5T+proTULei7qyb6hu1v0Y
si4ktTid29d9Jmpa/iNdLGYPUGQF92t8UW02vHw4fKqrePWiy+I8vdUtmIrnlC2yZKYKl4v6hX27
lJllFNujd0PT6/khJDMuPg9zXgQGqa1MHHeyHfLjdPP2lhMFn1omBhba/db61O/q3GaayaGFCoJm
854JKJPQWTxaGI25qohHMVCChL1lMOxe0zZOIJkbjTZUuuNQbHzCaAUQMMjb2UoTpfoRCKWndJr7
WBSwRpKdqeymwokgInp/d7lcSm5nCA4zqdZab80FmT8lXI8JaXcaBBowVV0kDKdGQiDSj76M+2Ac
efOYJirqD/NzH6Ba2cMs1Oh6e9AdpUdPAvx5lTNhiGpA6QlYKeDlb8mnemogDW96aDw/jRT+JFQw
hkMARQes7v5qZ7LG9K2Bf4qgp/PIg7G2kP0YVzkX4DpCyg7lBjMM2ER4bu67QyXwPrhF3BK711C9
eBwDuvbjLVv+siMvObt7cmHZbvkFyAYuW99sbIxQd/494KrgwZvYVBivTScpjN7PXyddqNtyCmbl
dVya2X8Vw6qSFrmSMXLFdEJ/Kvrh0T6aGrx+uN2XvPeU9W5HH+NpTX/AhnQduDvPx+G9TiVCr+Cq
z24D6mdTOhQHRoYbdV7PikhcPa7l8A/w4m4rcJKrSF28S1Lwk2R36cyYHrvwKuEPWrpUWYOk/Lur
K/8KcEgToIVLanisrZX7XYBCQI9y1cahhnC/Pajoi+lnviWTvxCtV/WNb52wI9K67Q+mcxGuZCD8
g7SL/6gWI/DVALEzezKMb06wb8AprqiOocmyfJAw6c7f90WElgcqBr68YeL7VoTY7m+SH84e3TyU
WgfXsC+t0y9Bsgqd+u5EBKuPRlrvBmRG7pF5EOq7QV3PNxESrgelKuAr1rCMWHVb1Q0F9yvDKGNX
7xhsd0XtK1Y5z7UI9Rmou8kYEoYHlfzRe6QFlMXJVaNP8FWPiCti5F1gz5+BRib1KB5EwbuE1u6g
t2hiCETS1IWw+pAtzE8KzG5N0zfXSyW/t7Ko6TqMdBAp8QXM7rU1XeBwnVlDxMmtUBg2ImkRgDMP
miEC3AE3ERNV1IHO0s+f4D9CNsFYNGBpBGuhDORXyc/sXnp78GcnB4ID3veHLcm8hCZ++8/v8jPz
u5hf7h7DUkHnsEYy0BRUcOOLNTGiigfx7BCZ6OFAWTp8LCSCMHAovnoXEygeg7NGmmu/Kz8pO5zU
hMgfDqWz6LhfKigM+9RaL42r2qU3MF8r4yB8dmY4PxUsGLBu4trmH9oagVE2i14mfywv5AUVHwyy
WKwnq2n5pOMsM7wjOwvJrpig/XR4zOEp//eXqpNyCJ2XsbQk9j2y+UnG/4FKJFCbewQPq2gPG3cJ
uG0R4VKLBn471rnU+G1ukbjZYWgjRSKeZY/MBz7Y7hDBLHDTZtKX/iBfayfNscQruHH56jjBMGvu
IQYvrdX44E9J/sDon3HXRRtM3z57I5IpEfRtXYYGFlQUQwj+FLRVGYZqdU588rE4JndyrvePTxhR
j3NhRFMPUeISTaIRjnWtaOUDd3UqcicLAiiaPMwt7r905QaOJSCzvtZ2V09PvaVWSuSf1me5tjaq
suYl/Ly7j/lDZpMZQysmBUzdLnZAmN9p2VeHqp492ZwdUBhpFX07hVNVj0AmqySC++xANDOX7Ce2
R24RaDVr7J42/zwW4e3hW0znc4ZaE27goN8oz3jmORFvX/qeNqICRBV+leCfh75RCRn2HC4UzNoO
gm/oDtDMUQ1dpTNlYsVgY8y9cCTFY98iALl/f4kspyG0VrtdvoQGSM7rWhmh0HvWJPiOOlG4pPD/
uv9gNmVxRcFZTTLpiFtnSGoSrMaA9Zs2yg4LI+TAfigvBZtTXhDRr9KMWYMUZHqL1IgT/60jmukD
jsQFUh49Wq8jfczrjGoSgaOQ1dttGa/U40E9iu1vrq+s05xy5Zkq9xb+mcqFbcou/5KcShyPz34L
RU3SvXPAkiu1AhfxTSPHrAkeYIsc7FEigIpLzYeW49e8Y8uRQOPJxsvSWfwdFo1Z/v0MFO3qb2JQ
eQ4SIkBZ5y8c9KoRA8DI4VHcRPO1saDG5d0bqLrWMSDmdUFaFsr8HCJWyu52yAp3a9eummWUtLJe
0GSDXrQaNJgvExbShwxUlTgqh1Tsj/jrrLTeQ8XXBSJQTwvmEqyLRMQfL4YhJS7n3HX1ZDrQZXJT
L4jO62oLW9SFuRIWOKuBKteiMSOwWKqD+akUR5LDvKkjgIIVE5cuzo3iNAYKqvUdNIAOLLjy/Uzn
2hErrHJ+C842pQYCSB6+3rscwagdodX1J5Q1s2B07k+mhLmUT4mExHnOn1C0LjCz7gWHXMFPbUz3
quzurYi5HcAjsE8iz0ZeAsPJgH4BjdA0jcL4YyrogklSnujzWNConlRaIoTcVLnymcIY5vGFgi+6
YW6NpDdFZCEVmyKghV55JJ6GmKFADTCa6nRCV5WUDTUzJl1OWTp08hALb+qYTRVLixrTZtvfgnBe
lbTWwpYstTnVc8YqWI9Ug/RZTFn7tGOymsAIDU4fr9pXFxPvM090RJkqbJH30EdqovIfbwkgh7sk
c/tvoRkCeFl9mhuWocl9dBPtMIb0V3hs+S7pi9i3CslGrKDJ3OMNsEftlP1kmmGxVf2/HjAhlsSq
XtJFtBbMKU6ta37/5JVygGmOCjKDwzkKvbOz+Po3bXQim7Z8LLOKsWzmQ0YLcyygU8dYETz6Uwzf
v/b8BaKM3fIcCDPO12WBAQSaxiG4HM7Z/zvEHXgLeYljYO4mDVUg/7/8AWFWOKbBXBi2eT0hmURS
39g5pFlqpy4eR1Nn3E512u2vYzpdtKc5NjkmYD9S2AxaFX8aV6wxdBD9F9ACfc5Bnww3CtCM4/5J
N10QECVaaOiVlcBXgjOS8tQZfJCIwheIZp9li/sxU0+YJImZbTOiLFHb+ei0MsOOnoXRxK6RCw4o
S8vCGFKstfunaiit8jMqqZCmoJLUi0+0daHbrQsgfJKw9s30AiVX4QhRqZq7CMwIW0WzOsNDHPMg
8RhBX8hQXQ9ZxgRpQ6er5tZLc831aAlpvAYxy07Bb7VrZnmwx5YECCHKToCb1KaBpcMqhg6PSjxg
XGxh7F8Iap1HnhokDjWGiFJGUB/VWMiSBmTDiv9fjvHmmSETsXpXTf5W+6RqBGcBtu0bzBcuy/U+
zETEiOqO+wpitm0o9h79DJKqd0NyeApDZ/ryZktiToTw0ivVMaf4sHoExu3qWdGxFvvcEqqxQznx
BOQZ44vdoWf5/9mufP6GbPLa4lwYBIvA3B7EaGCEvGx4dWJG/K7SZvWJuaLUJ/j6HvZ2Rj+DSPnP
ATlHl+b0JXIL/BrsWIc3exoAO8muDwVs5IPzDij18tUkebWPqCHr5ER9q0jMxoK9owPvjuq2JqJv
gu9vKLXWvhzN1ZBxrZUZXkTnVUE6e3G7XSe7Dx8kNKdLvc8bKsQT3vA0mu2kUW9vGTM4p5bKyQqb
JfMgOhxh3iq7EjQKDLmflBJQYvxYOBER8Wtuebgd5T17lIebSamlv/Ks7Hi21k66ediGLU8b4RxR
E2yUKx0eNwcGDvFycJtvLtaqOD6kPU2jEdXze/rAlKqXOKtASRS5YgcpmRzYWbLsc52HiLp9bwLA
LciscgzQQDOhEfLMkTu0HiL6eWJ07eLIJBEJpqEEj1+agKByJ4Z1yg8kJB+O6gMBLvJK4hZnfSku
SAXaUXwophXuA2T5/wVZ34hRXSZ8h3UeayaEN+by+9184UNzlAgFBO3xp0DRi/QMXPVT0tF+Dx2w
4hi7zJLJxMr2158ZIpkTAy2kDyKqhb8twTdux1v40zKaf4wUebAtwWs71UKYF3/9n/eJFR6Y2KiP
dvvqZrpvYnyb8bBjCbDKlEGVCzoVaGf+FwpsZwyx0jh3lRHt1EfNzknIcfkX3+FpEQ7Kkwwva+0k
h7PkkWMJ8nhxs55fINCyyiT8+DBBulOJDzcoTy2EYe3fmkDjgjO8L8KL3g42nKmd2l0qwYojHTM8
GtS76qi+KbI/wMACjLIdPqCXManKWZijiWqLLmH8x4I50atGfo/cOypF3oCuLtNeh5MewFMMnsBc
qCAhtpxKoVB+N/Mud1xSXLURWwFtKBhay3y6fzoRc5qFuwKJdf08NLduM8GdQW3O51NziehQQrip
dqrDNHP1z9qsl5EOGELX6h58EeAj9wJRGy4hdW2zfQIWPD4LDqVSslzMW928AsyL56sPM1NTFP/P
w99Zw4nWmG9ZFURj0hos3Y2oh6TLKXqRohWII6jLQGfsU7lvcd/OGRwxYcH/2AuqsL1/GOwrZXPd
DQSoxKl9HUcjsceujhQLgHnnHOKlm3kZUV0heafu63rIoWefdAVxVD9vtepUAk2wwFq3MQIauFBK
WQvgBFWO74fzaosIwjd7Ep5kgmuKTBO1zwgRcDOymVbGhB/tddBXFmxxOp2Cv8FB/LCXS2TEtqh3
1zRZxjCJz8tog6gMnG5/XivTMo5W/bLEm9rfu+q7K9mdkDdlocunhQf++Xrjy0AyJXJGNvXOduDH
joVTGPpZOratQu9jCIcQhCC7CRnl36SFhcE+wYV2kmfCQlR/pL4klCLLaPiBLzxZ8HkKOHRfAtA4
ijnEKvhr0uQQH4lt5GUyJ25DZYDh3IbmqSy8LSq5OVGTWwfYxxTYnYf5EtrJs9+yKIl1+m+2yMWn
tSJE70wv1Lu1KPu/Cn303A2iXJW9RmKdet3FIfYhQBpJ6e3nh2k1R0RJ6hTYMyBbxALTOf60Wr3H
vjuZC4sYpuZV6SF8o3fRa4mqhb7fiSDFhG9BEUOlblqtau6Mtp46/xDkVY0DulxVSSNIc8ccWsf8
+4bpnG1ZTqI+X7ZLvUGyTcUDYnWjfomgNva09vyxq+KIM8ukE65AyD2fuTr/5O6vxsYW2b2FE73g
KuU9y8xZIoTWpoIzehTuBcrm3XZgCh9BmA2Z+/RY3ScUqP5QclguvfOmGcVX6Re1Plbp9Nsoqgtq
xwaMvrcEm0OeQV/+LONhzDXmCRUK1fZCHxNBdT5f9Xaa+3pRlSkchTOrwjp1Tp0URfmDipCXRosG
iIPiisaCYG8DRxr0yfXtDt48ceRodygJvvo4PZwScbJgFMEKVYWvGW92RE2+KO4bWa8QtMp7vC89
BO8fL/gwcR1G7yJKwD657JA2wr87szlukLFQy+pAFGYSY/EwP4GVS9fEjozLCBRAq5mKYn2GwxXx
N4rqYj4FDNPTe1UeKugc26UQKqPTAac6E4Jh1yfw5mQoJ8+l9RunXxd9c2iuwZbPJ4yBAfyBguTb
wmVFtxJlSdpQ+9NDj3jX2ivKdeTT4SpeEb85oXcNKFVM6T+AI2jFu2zqWXx9bkP8YBV6biVhSy0y
3GOqMIO0OwSsULNQKG4RPjhWqHk4BYGne3+00/ocjGdGmJDDH1CU4Om1CtKf5PUp5LQ7Rmtgi/7N
2ZGDKVjlbgqZEF2NUAeaQvKQJmF8a+3eiI3feA5JD/TSKCPWiTNqi1ss7o5AJPVTpxryGkuH5jtR
lUVSyDFA6zxOiWSb/ncqDlzPR1xLuPg/G/zhGmK+1HYhv7YUmYA2t2/zr6/AK/YfER3ysRmf1CIf
O9xOJRFLpuV3W/BfbNspHTcNB7pwFktQPeBVLaom6HRl66VGtRjCGfc9LfuvsrPjJNJHaium7P2i
QVre9tsXkNlSMiKJoLZv/EMyM2WyTE0OZ63Z1u2/YwZ9h3kKNfyT/JG+BBmBCOgBaIkHEtB8hlhA
ulWwZTgvuy4SCLObt6MNeJooy1Q0fKaK9S7s7s8qpi5rNVKVrn8W5lffX0M+StZIu7Yh0F4yavl0
L1IA2P522Q+OQWhb6Q8ismwyhfIN6+fDA7fS9bU5GTo65N1yNs5kfKQfbKefAKiBkHnZWRnOTL8R
s58tZQ0+J5o2ptcWc2jR+cguj0htS7sP5PFCwQDFaDm8sC6JdC6w8bbKsEU/rvRJ08pTCAAroz8s
09+hNBhIW7MYmQUXNNjP9jUSNWhndVw1ZdkbEG17T/wZdEMP908h1ssvwR2HtLrJGVAJsHWjC6Sk
9GlikemOjNfLAh7JwXJ/7+P0yAPZICp7yBBN7lf0bGgM5SxtVihnXgLLfZOj8E8qpnUKGhqccRD2
cVAy7E6buOOUll5fspB/hPpp/kkLXJK8ccprzPDm3S+v++lAhDlBDrBWyKGF0EdWTdFP9f2FWUKR
nC1uDHDZDlRdvyMtVZbqcg81nyBrMX5YsdQ50I1acrKHdpD2xnF6E2ZXaYPg+sZiHwA5NxeysoD7
53LRo52qbpN+1uyIVFiZu70xuN9KH12irZbSi11+leqhDFWKfg6NfrGU19sRYOGHZVLuL883oTkw
SDdHbMVfBZzimF7KsapKA8sb44SNJtZxRYL41HwN0aTIwOsKieGyIoSUEYGMsThT0vty4ZwtZES0
+ERUi8CXKdZZBXBgYL/6Vo1RZh6qikN4u64gUBFQ7XADpNwvjm59v4GVIk8s7EvT7d436yCvE/ye
o+m4GcWpx4lIz2ddQGVRTe+ab5k1J63DqcZNYqBK9/r6tuO2Sx2JQolqEo9NJfDQFFDMKE49rOCt
MheEB2l4khdzhUtYaGos/e8zYRL7TKg1lojJWAG9Do4njmU1XOT5f8g84cz1Y1RzjcdGfUGfZ6vD
XDExWYexWXW05ptXzneFKgtndYIyF/ny9/O5lY4IvuRt6NWg8mk+8OGggLGNY0jsMng8y+/5EEEC
E4pI52R4hS5KOt5roZENWN6rBDMJemvpiNKSMNJO0fdhqIC69lXqWgslyujAzyCPJ/NJYi4jKhvC
tA9tF+HjAPMwdFh8xBEo60uX9n0EERpefFOwxXA4u0gS44I7EhssO04I4J5HqJnpdFNOpSKTEjdK
moXzKRYiqBPKqJaHqZDawNHPGRW1K9zCd9k4vIPbJFDOxsGnR2A0x0vAixiWCKYiullBr0Rz0/C7
tY9jDfhEwrkAbp/3SNfKA3Gc8wf6S9me0piUl7m3LHOOR/BPuJv2QwLzxllU2loiGrqJpULMRw7Y
/8XjrFQbygrHoz0m4aHHgNWmvnrmU9dC8d52l9hUNGZqhZ1nFkuiSganAVkXb2H5JLxfJh7pqtyV
rnhMlVEwWfIYkq/p0YnBFVqNrxla6Pk1TFd6EprIM66dQHR1G9REaUlM7oGlxXCi/Zt0l9WNUGyW
EttgQx1h8O4Zf8gm0M96g6avlRE8U1o2YPGz+nitedaI/m77enIKX9RQtA/e5AHszb+zm02os0mS
W803qLjMcvtUk6gczf0acLATSJa5Tbz/Yw1nij0L7dkPwGf5x0XFsjTei3IWaC7Hk4NVQsW/BaSY
G1hS5P6YxprXAdjye2P2Mhh3njH10RD24QMiOH9Gnx+c/TV5PB9phlwsaBWebmNywGAGFwGXU5c6
s7NANb8sGCu8Cbi+8GrIDcKYiu0VC5P6oD6u0I4DL8zKtozbbI1e1P6d0JXIiLuuYjmfJ946I7TK
zNBa75h2NtrE6uIU8Jd7ABpZ6murYCq2JtQhNvCB3HH9J9zU/yAUUsLclgGHSZureQ+F0YZtRN25
+Js/GEKSSeP6UrYj+FNjGUeTlC+vnET4YZu7NENQsED5pR8DiRs+yl2wcaRO3lJ+COXCBabSETmM
4fxlBa8ACIm9J+MqcKIozsufb8I94c0LZKmC9QkXMm0EhE1CAipVIrFlcOjXjVv2VAQAf32weD1x
gELxZ48rYB7oYuaWuiK2hKKLYjHzTJz6KvT8zDn2/53LMOzflLGQUSxyJcTvcNlVxdCbH0wIzw9k
j8OoqHeIsi6BN8DZuBN8ehA1qobMm7/+VYDXuNZ3Jk95M0h0qwwukXQmGs5AnkUiGAiU1QNGuTUT
EOs/p814VifjLymoJO20O+PkpSS6uvauk3Mwfn1Iok0kGenc/UdHHRTBwVAEzBcbUTlhW35DsPFe
F/dgiv8S2cKlv71R9FyVGAplu4q5y2r95oZTm/TJGgJeQda7IKQGbNOxJbDJIYPaRT3jOXK0BE12
GcUN2unnvJ3j3VfhNYte4JN+ki9JcuPsfepvptl4jUlhWvw5mB+7PVLC89mX/juOUyCbm7E1/fAi
hDVPIl/E7AVyzQEgpQylenuboQ8JnkGefFAQeuLo/AyiDF85gYzyJ6Yww5abw0fLEtpfCZh6f7Nw
phUdZ5bTFx0v+12ZgDVyYQFTt3daY5V/+ADzGFx98bIcEl3v6x/M/kRrzoKaWGgroiiXdH6cmDbi
yo7K7q8klaSUVr3slaj1GEO+0cmtJ2eVaeoWkepHck/qNd9h4Gswify0hiQFo0TQtmP6+uqZn9eF
osJSD9ZgJ3o9PYk0X2RRiEecB3ZnCAyeBIv8KMIeA1U4nptdaLKwsnjv1Oa86m7jugueaVnzFhS8
oPT62rU2ecV9IL194PPJJAWfn88pyefibz6HW8zh4cTJsy/r0FBDYwpPoiR0yAxm/sCCdP18yFSt
vPJF+7KiG3PE3Kfe07agKbV7NY+Kz8cTE9EuFkmcQ/ucay0y0qjYUlxy27F6Z3PtZFDkgMIGWInh
9PsO4pD7b2oMDjge7lW9BDVB4mb3wXqmp1//sxIRpa/HRAfm2KvWWVKhiiLi5cdcsGEmbpa41Xvk
OVDUze4rEJHWxpRGBzw28H9HCXf+bMv+FhP+MoJrA5SRAWZMPs/FirkRbYks3ocx61vT2OkpLoaX
o6VR8geYxzqZhPux/2SToNJWj5+BEWu2i6LD4CBQrTTl9vvdOryzseJPtoLxH2NULzB8eQGuEsNm
6ioeJuUH8MSwDG4rpTYxbACKnfpx4nEHZf9k7+0Qz68QmTPq7PHKnSszVZJdzWkVhZr1DXAXgnOD
5LShelsWogSM3x8CqF2b8yn0qSCLFe80Vr0KL2LKBh3sVObp/DVPu5Q+CeYEd/tcYlRp7kIq/o/1
rgTfjfJSgN1mjjyYkNTplIoxRse3/qQf3prrRGpm0nwpfn6Z0Syu2JZStWromjF3lazqzXrA7LiH
HAkw/VqTCE//HSwAPyfYRHyIh5gtqlGziHTfazs1+D1gDZac/JxcUlHN5shDGtpbtYF7x+lyqqzE
Y/xJy1olzsejU7lzTK6Taq80uFY2lzYus5Z/O3PlLHZgCxJAcJJheX3vvGaVGqL/qMmTbFiGiYE2
IQm/Uj1sJe/C1AIgoj5189qHP+kFFwQTlBqd4T3pqvSZEfRFjvaZgsU6mzstgt3MsQQwM/NLghcR
1zxrcqyxw4lttzoj0oxzh2X8wJA9qwM7mnkKTaqFGQKuXUfu6ipPEIgHx33VjbRQR9j+oHaZ7xIJ
IjxgV8dS1yh7HTFMCQevmOtcI5S+oPPN+eGCsfnNktjYXO2qKEKG90pAt3KviSrJ5t5GeZ1ZSvCJ
AZPuzBcDQwaei8Rcl0gZPi3y/O+M6hZT9d72NdyHemXTu2HTQbBk5pvF++6ZSdpl/cGB4FiViY7R
8VcIN08J9IdWICPQxtZh8K0zAqmFU0imBFprU74j3Yv9ZPfvBq+/NUUUPT0Ka0DjfeU37CY3n03F
VKgVlHc3WbPUNOl7VWCXGuEqfAa5hFigV0a6Ih7Wt51N6tBK4BcAfwTws4aeEjCniGimP70gcw4R
g0kY5m7VzIa1EEOSgjD5AUaoLaiUs6HPGX1Ba/IOf5562KP/JZ9P6ek+jdk6dGS5BDluKfzRVWv0
j+O89b1LHTRDao9DEYYp60RB8F+y3aYFnhozaEAUAuzXNI6S6vOAQHb2elSHKGHUrRKk+VF5TCZ3
XC8RyEsR96LRPZFPFbkn8H3lZHTi+gwxaBudmZ/fzeZrEzyFIFT2gO3c8xCrik2vuzPBfpDwZKDB
k9PA/9Ufl1nKDAKAti6i9fuBrIe9uiT/zLcwQNucYGwOOZ49a5df3XUiWPvvwRdkC05R+6VBCX4j
2350syVT62mnUTDtMBMU+T4owMTKjaRqRI/ZqD+SXup6fcpHcsijQjSz3E05hLPyiF+4WF7VDvPs
Tnu3RBTAkBGfW2mRudDqfat9or7nfjHMY7d0dmqPbEePCmuY4ETjdtwPSLkDBvAODEX8KRjizQ2m
dXOhfLy8ZFgPaA0ZZDJxVu+Ydb3zpKVhfEWqGSS39bGjn+LEhCsRTnYLQzOv9eoQPtTWqkYSnfPU
Ez20yP0DrMJ4LFOBJfckjXsLlRbH0rN/DbNyxHf2tWdVrpuCnM5F375B5IlFRqrtVbTuzr/xQ/ip
XYK8iPsj2omNAfrpbKlS4HN/ohcaZNfKZ3hEqc0DskME/7Mkj6oSaQgJTdlkyD/ns1uBpLjUw9CC
pt2L8qTEXupNppH2CW5VITK16xM0BCbLVPGMnZ41adlPTJEAJPevco97BwioGbYEU3SXtZok06yE
QGgozQLi4QRDAiZDg8jadYEUMm0k4BzqpZc37bf0/3KZdDOLveOLrHvFCBA5ctMsdDBFwxA9Vqrv
iL0wFLcBGpLvzg/KTlGgU/n5fbnxLuky+CA2IYyqTp/uUouDEn1kQhPYsXtgBMxyqLlLjeVDl5jf
qo2vcha3dSVfxRkM98UnpGt4d/VQ3QJd4/Os5rkg0lPlLkwu+nDgUQ7pXjQRH6WqmJ9Xci+5Eq66
HspUY48s8wy1GVprzVljkqIPuTI1gXJiUdxT9D55n21D2219zPTzMKTf6NGCJGVTRkHFkamFowSn
x6Nz9kYJF7bkLVUFHRVoYQaleWZnh4i8ZE0NJftXZm6+bhMwQRa1UKiFT0G0NKYiO3reuAfZlzkH
RFhlJgUoDQsaMDva04vCFF5a2t2YM9B80ilzdVQvuLLYJMtCYUoIZ53rCUVBIPY4YI+Gpr1xuWkO
b7NQbX4miinH35jKw0yHdsDNBCWxTwr2+DxWkjKKRKKF/jGBEx7J3qGOIdwsubelKCrCc7vtZi+8
Js11gdt6MTnmJIlScVxHcJihkrXvas/QeDvjw7sFveLh8myWpbvVTEc7fIjjPcW0VvI/FlqBZwl3
PpYoT7MpdGPy6/xerRabzsFfryoh3KZn0LrnJopbWjUm58iFphN6pyv4fYDsk+CqJYmSP5i+tMY3
hR+j7tMuDLCMjzipyFXZ9JKEhcVVlRwi+BKP8lRiobrPuNKJI7iIs+TK3VvbQFlPURA5gkCekA6i
2I85JwY532ZoB3Saaj471+V0ThsoePInhUiMqH6kpW8GKMQtigE4MIB0+0yc1qWKD9ay52lSugTt
cXkgAOxPSCIcTL+2dNslF0v7DXtR8W83sL64DYWy7uFjCLJI5mOb8Eg+W7GRYmu7oqE39KQMvDON
5rk6fnI7BCtIIeL3cp7/4PcPJ5cV1MgKhniRuQfkEvU0iLoF/NxQzKA5SaipRrezILaEA+/KwM3L
uukFqMdN9yPoKqX5EVWUHSy2vFsirAIJj5o3YR58s3AyfwtZM5g1oeyQ2yodC4vbO9FC+7v4Law7
NfjPwblHPHvXqxrowUD4NRTL8bJznfYukNyuB9yqWPxcPfmFhx1vt5KYHSoz/CaloMS5+HwjKoLT
K6fGIHeEEahATi/8maxMlajgsBny7knJIEZzOMpCwZR18zGKWRMDMpDUQiDdOWhpedS3Dycz3Lac
sCA7Sr7Jc0huBSuacl0lgkOs0YouCxP4TZ42N//2QBQzWbunSeWwpCJEAiyxrIZbnZVcUiXHJ+Bf
ZO3ZOFVeXeji10SS+s4N8vovc1JJEMoUl9PbwjGMHeBFrD4N3AGwR2l2m0HX5r0zAX6xGjM5Gxc0
Hdc/ce3C/Guo5Z6x3ofwgXQ6839iPqUKMyPIAQDrD6SGSxcxAmWR+AAE1xFjVkRciV5JJ0YNx7zf
vy4OaLce+kwIT7WFJ4clgq2Bi72JAD/Vzy3kK8PrpWjdh43KR2HgHKXvgsvt3IFhV6/xYmCjOUXl
emWp/lqSRNl6yvYKMPHUVtPs3Pbgk3ijCQulh2PZjStRfKYgcdWNG2X1f2F8suj5u1CbIQYEsBgM
eAq7KyrrPNK5Xg44CWkIkm4DmNWauIlhQgswug0LyRfNmONfbPBASeJttwk0zhgt2ARE+g/wpDga
2ReJ/QVNJzA9b7YKiYajP05kzO25Fl8RdaE7Ws3saC9map2VFtMVqiKs8DCxPZI8jF2iZ/MpOs2C
e3GX1XDwjmdN+nC3OFAGiCg7/1i+buyXEYkprjNE+tkyQU3usvAD7MLdl1uNXAqSeW4RKMx/QstE
t+89DEj2X7JzjPEPaWNpZF6htHomFKl2hACbnrBgb4Ju4z50tROw1EQIvHsadEHbEI4IE5xwfrSq
knkvjUcOoi5lUcwy5vAi7oepfmmEtOEKXPARt2nFvdMsUukOLGfd2/yl4K1uQBuc34H25d/oP0gO
2FPD0vl5npx0FqjrrgtQWKE7P+29uHCNPcItYbfRekzsFfG2YMG7zk7JkcWl3gpBgqf1nS1AWssp
f91IWWm/O88sPSNzezLv3yennNiQBtExcf0mm1R3gBZtLZJdsCfBHNEmjYLG3wsN2/3NiMy7K3uT
SGlQQ2qDDSQCIBbPZdcAbTkkQCtEP4e+bj0UOPwfa9fWnWWoD8XPDnK/gGvA4QbPoRjrROnn1Rp3
FotFd/U6MYl8kfulOArm8YxJT/PXY8TGWbLL4yiQe1M80UZZl6fEcnJ3pYyQAG6NGNQfIj78x/oO
TbYv1AvQDQR2Z2khFdeJmm+rNoUS1KzCOak8gxMOMP81c4svXHYp75nlAdtrbMnBfR1lED0XU6WJ
Uoo8Y5Ac7HymwkEkVtcIkDCq/idFkX0F3mheVD8P3lc62l5Jt86NJ4pvSMuOLdA16Clw01wrq/Mv
gE1A3vSXv3eNqjX6Vu3ea7hwpDv4dt7I55ROppc1MaLklAuUA5hTer1MxtOFJ06u8oVxxrceQ6Vt
fOZZ0tKHBJRlLNjdUBpYBv2G6yQOGIuhaySbfsfPLOGtpfoQ4qQj7JMyyVp4gPnuvAqKACDONynq
pqSOYaAmQQ6Pb3BgqPKFCVujangUTgQRGNiKqzPgQHzeYmlX8IQMkkJTpTRwt4xvhRVheuSz7ob3
pMsa2GR+RyzG06EGjJJCECRSqBqOJMGsYBH8vdVu5A7XpSsqbMyzU0mjsDNK8ERddRqXhzJHKj9N
VTvNFadh07YtlvphosXIVixF76uiEcAOyum970RX1RCFTKtax1VcN5p4UDjRlBPDR4KKD0jKnqh7
JX7x+iaN+V2JQtAKSzfENNbO4GDVbcyNc7Xyl73NBQyvzFculvllH+eKHajC6mF8r35AMdZ7zmaa
NOjBAawDRdyHqw+zwy1SniC3sMBGAnXgklN/ZQIijhhbst6CODlNm03UILkIrzyta/uKbgmlpTbJ
VarocpDc2koV4XHHUl7b7uXB2co40KsXv0baYSmbhAQdrNTW5Z576VbPMhbRdFodfxSObyaswg3w
xg7TbGItbHw+Eo9lk7mvdqz8eE89zEry4/m+BI6c2ntF1CYtZ8K1Zaj9Gmi/+QWhh4zuT/K9QAvm
1VBHscJ9CUNWxHudPxSvTr3ZaBXPiKeS8II7bXqdDV21xnTYEORqz9LcbPJ27ituMTYeXI3SCPFI
Yv1ANevLiTwo2ouT/v7eSNoRBtC8RKWL56wtHJvc7fY+K24q77H09Weir2pboj8EeQtwv83yPK/l
6lPn8RLUI7o+6vyvz4WMKGpnlidamc5u/v16yxd9t8gIAqLv5fN4SI1jfp59gRa7QQmIbj8a2MYE
IIccj+5tRpPIMYW3q/TdC44RpbtEjdOTdp7nZGWrbhsR3u+j423o24lvjRFTLw97GEXOS8tUpW7q
BUj0jWG9biVr2WLAiQm9CbuuBdJxqDvZWTVJgNY82wqXnr5XzrtVqdDF/F6t05h+IHfnIB1nF1xE
FsgNgi7jo/ldiPQrsMR4/CO7GMcnmHnA2lrhQgKPevaMMX4E7Iy2vpPY9T0xuKyEyf6VnvZsqvyj
L6e53UVW+XZ9dpy/oS0TNqvHEQSRTMpVUr9pSb3oEcexClYCCm16ik/as90GsWRkK+1Fkf+MrSXX
tTRd0fUHY4AsvRlKnVnCA30Ka8sBFCPzLneDf0jEFrMqRFQOagd/C97tVYaj196NNDVIGjqm+jQ9
hgswklyQAKzBlyI+sRXTNpgLEhVKrne4wH4gMRo9wybbKhmwi9p6i074KXdrp8DGR+InDa1NYDki
7Lup0NNRqwk6FfmEd6ASLzHgTVGTXgIzBJp8jHwgu99ZdaGbMnot9JAaDpyV+jEKBaHjF4uCjayy
Iywljsb2gVEcxUltdjy/QOCA4t4AZp66/bsllgZL8m/gB4Nzu1HQKsomkdJDQNZXZrRuc/jrjf2o
0Ak3qcuhJxAgUfDr+DaTzuMGCU7JyuxyM2krvK8YRWN2EtEQydPrC/NYdA3iZ4q6ftWhORbfSY4P
sCvXMgBHvipthWnFZ/SNihBKJKtmuf35ofVyrKfYnvRiEsCC5uxMiLrUdhnq4EQfHmj0pKn3dtEW
HNO6Lz4D3KOXWvMx7kQeHauxzZnoVzokHggvIHBpCBu5ZlZ8s2im1xUuRqSlimzi/iOC5Ci0lzTl
ydJANGaax1cgdopcRvuDmQ+TbppVkVjB9FWUI1uepJ7h16qAy6a115MLBF5oVsnvdirPAUiZ/ZTD
vMOntqlqyioDpjMITNab6GuHrc7GEfrrvdq4eEQp0yDkHekNjmACjdzgNfNvGWCqrRH0bo4ha44W
UBdRneuoeyxlDaxhKuPCLQrmghr37nDJFMNG7hhAdbZcGEkmg3/JP7paH9CL8/hQKsfJTv0bOzru
oaBe7eV3XE1CZimNHhvfeS+/0CyIp27YqHcOSii8VHw/nKQXMJMuwpKrtUeN9e+I3Kn99vAevVeh
TWGIlv6pwV7kS4dr4ced4FzNm64i1lxwlR1DzBhEFkI50gFflhpUHnMlwq6xqBx+ynDwOr6UR2NQ
Vz5AhhzPw5dN0p43FQpUJm+ogkRe1TdwVunRhsrbluEN6/3GGn/jFXDrhieWm/K74+3uAY1lCpuI
qIzecmJSXIuaThPnUImPZuXRsP7Dqe2yfmgbJiVKdsWBOj6dP1pB8+ajBDjzcF1T3CatqIK85VBW
/oDaC0mWuZUU4RIzRFO18XZYRiMwpdQg+GIkt5YdEVcAmP0F1n46fBDXtuI61ocSykwDpg4K8XI1
DYPpCv23CH/EVjyC1t4tQbomebm5xXA8Noo0UjstD+7nilwqam/EAYawkxJfzS1pku8rSrUlzSdf
VK1jn/nnuxn9H12zsfJ4BJWj5oEKwlODndccpARUKQYUrj9bvw+vcESGnZjnFXfQ5rxNGiXlXq/H
6z8m5gp76VAKEzoSOasn3V/Jw947tL2NhbWXNHQfH/ndNET6wKALIr52xWxhjFcVHHMR6IjvZBFv
u/CyiFKZQvK7LztjPytgRQjE7TYbuWHqVLq9k6++qVJ+CzX2t6t3TOEJ9nC1vrKiWW/PS8NcjMXX
mArnY+L+no7L0/4SVJorJVV9FjNzO4YZLSx3tDx+qXF52TZBN8p0BGzZUGi7bQ6u+rmVJuW8C3jP
5mL0dkj6FnVIFLb0hx4jWl6qlzlGiPpD8zFzjCGEBt9WPi7SGohdeUoZgx6rEKjxepqHtqvu39Ov
YkcLLboFH/AybeJG22Y/Ee9kRIKxTK0XxblOiwTQoiv6FVHUkCJ9demV8HS0EoAdPzOLD7swxwW5
nFYduJyNXGfs6wkZznxgAXnzyMVnOKC0bcQLOjyigXVm6bw9nU5xzhJn8Jnul5/EoQ6CM3Jm2USZ
p699/6qM2znwatNJvLPfQWCEOZ3h8Z/daNq8uO+IG0bkWY5XeXLOpvosSI8/dtRpEREooEHCOsfb
wl/TcaCtL9sVqx0kzaJyR2xnnKhb4ftnThbPJDJuC8R+oDMvvq+ovgBngMNQN+st96TBJCvJJcmH
OIKfp93Sc8JQZpz5f/h04xCDuIltcQl+ghnXDr75CY9EuSkWs+ui7n9hCdHO1UH77AEhrnMHie2o
+9S98EzizxUOQEya/m0INH/n52+RYCU+7rcwJCp3z5bzVpkhOjFur4oISVw98GHav/oDIqhfvpwR
9FIJImSXIFNFqmvW4UCFjuywXy/pT2SWLeQNHUtOfEhDEu2qtysXqpRoc/cX3pjK+CbHF/56ExQs
OQWJgoR2Ny8KuD7ev8Nus2PmnU1hLJr1rDe0ekg6EKmXe8yGHNg2hTF11tcevRILdEOUSlS+vGCh
vgFev9xXDkhgPRnnMH/CIWdg9lJzOjkM3BWj2PAcRWqT0qQpQ+iMiDZHaynF6s60LH55toLpza0C
5HeBdl7MR6aKfLta/3XRq4/QHEXuswkC28eK7VpeGYX3URI8oMfd7/H4ZdrrvPjKn9LNfoebfYKi
Khr38fthjSMMuu0D/l9yiHyT29jnshOpPIGtkRHOaqw1Nnv3Ih621X4fnq7UEnjAxHfxnQ5rH3S6
hXLmxg2Lbj0kvtIi/qpWiWXmEg9QiGw7mX8ePJ6W2NUoBF/ymZhhY4RAriRZvorseMBKX7eWgQNv
UlA0aVDuInfu/mVJ0QR41CYV//qmfOiWnnWaZTMroKkPeqeFx4ceSWO+DN4f7++nvluhkyzVtMGn
nQYgpNzHuysJqT8yxIQkDMIB/sytp26pvMv3x6JyLokGVGCgNRB24zseRxZkbluPZfb7hT7BGrjE
zGH2Th5KDxt3O6qKRfrlIL3rNCc7WXUgjvk5Ds2ZFFUmWvvKpr0C785fZvXrR/gg4kWFaGyyQEUz
wqW8F3UTS9FApDhKz+DZkViknWlmaUYWqmwxZk0mbx01NUIhrTEchD9Z4aJg5nfH7mOhip4NAtQD
gFMDzUF6+8/iPp0XupDZpxu8s2STdh5z3zSgwExdEBrxAA0UNXK+3Zcrh6N6PvttYeaQ1F6DHYb5
8voItcQ4yNz02wmjOAD0mVCF0KWiM1Hc/byhLHDHHaIXeFgO9WKf83K5ByO6ZpKMlrjC8CB9wisl
1sOIzFJYZRQcVwkbmmCudI+BhVF1L+Qq7Omah4KzMXwh5Aigm6pCwVCe3NLKLktm6GvK6C9/OReb
WbaVCzDudHqs5PE3r0U6yl8aw7E2TbCEOFWszmG6JM1IWajGb8w6phejU85aoOncA5ZqFV49s921
8nANlQJAFhYGTyH2/3TDBgiITU89cWmAtrekwOxMbtC11n3rM4SHcv4mr2BwuJujlYDdwnfTZG5S
io1ktyl7CCc0H4Z1g1Fy4p09lmt1oL1Fh5HIOgt1QLoQCTDxiKyucwO6wmNImnxW0IE+Tj2PQkzM
rAGK8wKAHtxShHzLwIUPU+/kFC9P1N0UO3Io97hFCV7HKZVhWtNi+MIZF6e4bNg7IOndTeKBBkX6
QUNcwKY7r+QqvnDrNSfA90v3qIzDLuBfwssyQerdct2Z4iNxJBpqIqC6seJ8po2X9ptIkvBZd68w
tKfr7f5KziYUx/IQ9dQ74e1XoNDfSJzwRqJ2BhSH3xLlU5DU+UtJxb+RV0oG8FoiBvOXrd/kqmEy
N4CIN9dKKI4DpFVd1YUg/WarxLGYqJknFrQfhP7qyIIkC8PjjgvhLJfp5dY+PFO9s73UQ+r8ctOg
BRhSL+kp/BEiH4vG3JtzMx56ML9VLXRBJHCBtFstC0DqJdVyFuLVR38/L5RJBxP6AMvNBt3DN9Ss
/opGU7HBDeoduGPoUDRTCVbXac9DT4JuCnAy+Oso1BI1GvgXTlweW6KrXG7cqpuIngCESdQBYysI
Jhl/C1svZ0zMKGbk8/pG7ZX60R01K55cP+PRbvxFME3hQ1/fNDANVGgnOKIaA9EtP4FrUwuk06zl
5z6VdyqRvY7rBpVQ9SrWiHWDhh8rOHsZbXjjBzwCo1h6MoDWnHY/nehOIwAgHS+mdom7gP3wXazO
SuETUP2IOyGp/q7NXMFtlq9Sihh0RgSdwwqdNStk8gqk8pcs+UQYZt+/xSivbHfyAshkHuFztQzv
UGZEtoEIJdmZ1Sh5n+ddSqsxyDG86yqf1gHxlKMGin1VRyERUXLzsAuop1CdnWU/ky831H8B/Nd4
ZZbReaB4/0Q9QHNh+vbx49lgEfIrpwoTNZp5Za3w6miJ5RR0YfgmYBXv2xq+L0aHUM0piaF2TAx4
4+si5O2OuV8cISjz1nBMsGrKBcfWSgQ/xe2tTp61Nj4IlOWWpHrbXivrkfvGxxVCliIO2NKk3Kpe
HfuKYnlhe2x5OL/GpG10kKUUkNngYGvJbxlDSFv893SN+Py3Ld1M4G5uGpNZmtFUcB/deLEccMkv
Ykpde9e3lJTNggJft9s3SUUIQYTUkUNyzx/Z0gybf8T4GH3n5yYwmlU9XfFot08/vSCGUJZIImVD
FfEMX02YcsntyjPAwscQnWrgs09ASscDOA34/320A3lEL0xFzNZEx7J8hDWqGIz5sXVOpkoVYEdD
f+IcAl7RaUQ6Ax1DGX0p2mP9+o+1BAfSFnRrz7NgKtRCn+4mb29t0yPZdQrO6oHt//gVYAEuzgyY
ahZ5ZkJKu19ZCzjoxRzh7IJxA3f5HWedrcJ02sKyWvysyH5z4kBDLd+uTzbNL2VmUhjsrmelgccb
jrd69/ajXnJ16q8zEC/K49WmsJPinNjVWGsMvJeuiFbghlj3mx8R0+m5ArH+hHsxuGaco+mlop58
rvPWqF2oMg/vzx5jbb5eGVmIK33Xakcxuy22TogboqlN2jmK4UkguCogXot7NGaew2/dPui4HOSi
PnsEk8QIzr7DQi2esqBsnDY8Z0B6Vp0ct1jhbW8oSoNX1Zj8iGTKMbeA5L0LND6DVlbpz3p9hobS
UoHhE1vmNbtOZtqYkOHj+LiRXPoy7ZB/lms6l1eCaFFjVSVRenmor6uQjvYMcYl2mOzZaJzy0AS+
BH9GZzu6OC1U1Chu/sz9B0YSuzKBLrtYMJboRnGudOtN6IYurb2mbW/2oWPDB8W2vp8gCkpjk1V+
K2nB10ubCU6Lt2QQn+3U2a/PODlSFZGBWc89sL/yQXC6cUaqJswaOnoP//rwtOX1MGeaTWJoGg9v
l/1OrtWo7yCLjGVQjpdrx+kNriV0BpQRaJsQe8eAXd7w/3UUmYEE52wBY65mH4HUehwVu+JOYUQZ
X6ri8jGNgLhc6tuhGf/gtXChSeY/FWz8atnznpgrfYCkfcGAOf1KZMTBkMADSN9k9EmqnTitCY05
5WRc3T79Ctjn/g8YPiDBIJB4FJmGQZ1CIGHfAxPcpINJ2lXGRqIfoCgWk1OKj9Fzg53wVnN/cJor
94zh0vxoHtCHmnqxqcetCDdGfqQA0Kwh/6ndGFzKIhCGS/efOVcmGNiINhmbkHmZloz4hHHdWeWI
Xhqzl/QsIqs+e5QBQFMAIEFICrM7nudoJRi3wZ2D/wsWvxGGjRCfBXCV644JOtSVY7lNl7DJwWcI
dIWpD8hD6p0tjPuBHu96bimuXWn7sqr+NDPp1mU+blZg1dcOKUW2pINl2yH7cfro+gl05iZZLEY5
pnf8dvrJpBgvp1dFciboV/qyPhk1wIPNUriAtPhW0RLOcpzlDxSddt070+lZTEBo156LVGGnXl5S
b069Bm8KoegdgJLcg7aOYs1ISMyqBqMN0HZS8tpKrm9YJ9CF3AeBaOaAnb8K3sq0phta8jhIrtzO
ogltI2rknMiveBb8GbmikoM+3x4Y+LLzpjfYjvFyYrShjK0Z5Z+BwM1il906NcBzmG5tMAsJ386/
sKum2lHZ6NmFwgGidPIdIQpIi+Mn/RA5D/u2kxZ6F43neqpzyTaVv9yV63bL43e2MZeuEXeDrGhA
9kEydME2383c0dCTwjLQi+0mtclMdAJDTGAQwr+vBOd2sRTJHjeAuhEM2sNxBENbByGRy6airzzW
gijSQ5KGzojy+CxxeFT4uK4LzQKmSPGUfBbt/MYuuGwAulEg7co/Lju9FS2xYGY2m5C19O+OBj/B
4B2EA+oBYmvRIvD757AknQ5eHEdtD6C0LQHbEFrQ3T3JSz/MhC+a9NvU4vv3FhMnVMY6nxJiJL+7
FgXvKaLpOZigQpx9ahX/rvX7mNVgHmBIfPZp9zE0m6qfhLeJ3O7qJXygZWmyy6maGhHZR3RN0VAM
n7flzvEANEk/8ksj7T57Cegu4w0xzr7uSr0zagspgNPphtfC1dNBbBVU9hdmwxFdQO6LqQABY3kk
gvoruPXZoaFMjZ93LedYGq7I9RVTGpgpj9EaFGkE/y7QspOyTuDa8Y4qnepq2RyBvSKJVi2S8DpA
D4b6AayazjfIHex0z3hwpbSI7pk65jnD8W8kaX6dvN7U0MWEPt0++vhboRzHYrfdEP9z5nGWN9sI
sDbDPCR4X1jZIdQ4tUPo0H3l8/Kg5mVePXWh/egtKfnasRBZHNPkKg2Iezzkv+9ptAotRfrX14LO
yRWLcWkggR9zYRg6w9ZJ53IpXNgJ33Ze1Zj3XwA9Wuvojt84A7ZPjNsnRxraonzdTgwyJ6vwFw9Y
TYuG9gHEIj4NyPowuUc3aKj5k81/CC4H09UQCXNCFE06UW6BZJRdFM9/dF2+ZWC794dfOaezOgwq
WYXFRy/Raw5QpbMUnpiWw92lKRQIG7ml5ZcVMp2oJxf/oxC5KUY75Yq+BvyzVvluCOlp4T89ltgz
1VyffO9iV49azbYl1UIJ8KBoXotWlCALB2uwGIj39QG5gvFY6RbIfm2m9OzLyQV37jRu6TzG0M8H
WX5AKTFsql6gj0REbbY9ObEETup3DIaKmE1M95OrIzPiG24vPE033U0/13wW421dOU3Lr/PS7+J1
itPB30Oz+Ku//WV8gxhIj+l/m53o9ozDE/uU4ZtgXt3aNppaL4Ec4bmRnv9WX1CKDLxbHh9hAjF1
nnDmGdlC0VghNLIOFYMfgwuVZQJJ1Ns+GYcmD3kewFAH0qGnYpPzZ9KlTTVTLyX615HIpiItInBh
nlSjavjlaYdb0mCTxDn0wrsm984poqrIYuZMZE4IevKzStXCNWMbHPGZxxRYoQOQG8jlUD/+2ZJj
Yt4M95GAGPAwOwJqITxR6rMozH0eo3mTwu4AYHv/mB1k37KDCWkCzHevENeJdVUnsGE3PvJUeAWl
jfzV71TlGfSZGoebupdrh8cWcsVE1+knZfckizVH6pIueFLlGKitY9pxN++Q4uk2pjHjNfm5i+8r
s3Q5FS/nQqrhGCoc85FyA7RsPwzI5ekDQAVOI+/mo+jzBLmYWm97uRYw+N/zy3D4J4DqnVntyOL8
QEnpL+90/XmWhnNylmWuY2BJ8zx4ou9DKbVaK0h1p5zcQFp+nucd32/glucu7HVKcylE8qzaCH0f
BjZ3v1otKJcob1DOPsxELTUguJD57maoyooSxPiKDgMuYAo1CIXml7wdErLV4/gi5PwtkE/we4so
nkmDFHL4F+fM/QWoBDeV+vCo/wVgb31FsKrOYSqkDnDGmGOW1aEcAMJeQzstsNrU0NIh2caGPdxF
AZwOJ+t+Ud8RzqWhgC16/3SSZrD6PR0I6SM7lJgzZYyYJimJRgP0JGjc3Lh5bAtzVd2sorIRyEc0
/Hct9bKZFeeMrscvJE+n0YdHDNTnpiZYQWAyYAWMKfROML7IFroBdz/1cFW29iRinMOvblYHugQo
SkCsgkT5vmqmGp0ztUWTlbCptKcNprhAXS+OZMBnaQkecBiV/kTSWjLydAt8yWJuNTsUVY1lGS7T
4ywHe0daF5kyNJgrPw2ZCUWvm2cbCy+9Ee0G0D+HpjZ4xn01e+00WYs0rySdCiTXib04QK6hIgnn
Uv+Jy/lIRoXPxokXJCsv2auuFy2X4GNGltL8jkrQArb7NbHSacqrcFq8NVEnb2MODOy01aNSYxG5
2seXEsjYYPldJDOpt72mGjFlp9HAHpJEljpnCotpk/2kt/mrusf+GrOREEutA+NB+zOlA5EkxyNR
oN8+k/urbOrcGuqaFZqCTrKDuS7aIvt+pW6w+dJSkIB4VAY6b0Lo+gYDs6i4s07f2zSNXsH3Wmnd
2Tq88CZ+LFQXlVA0UUuN9+XbagOY57zk1/XA7t/nah57TQ6EhBgU/r/U0N0uljTvv7ahWERaMhNm
cpeboBHmZ9R3bYNgV3Ar4G4iDYplDldPCLoRwIOqbgRLOoRvH9s0WjB2z/AVzt/XR+mD9ux89ff7
TLRxaiE0F5KhCvi9U5sr+sO3Hpt8s5hGGOhDYwVnnRjleNbt9NP6jlEF9G811Lr+MU4FSLg8aXTY
F/OGs5MGJIDB4sTrRQ3qxpwkCmiCn6GJtptEEep/Gnt0hqE4PCbddD6QcahXD03dLpUkltQ83fLk
8PbJ/OIm6hecEgF/L7t/wARaKBId2yYn4jyMqV0B5CqaJUynoquIW0MA8ZyU1dYD1qX1ocLtHajR
b+u6tqJ0UnaX6IFqjYPotdIHo90kUpn+Z0lIGN7tEuYt987qtiyL6cOzTv6u9QKwG57dlxi5h/YC
eIBUsR3kQh78bsIIZiu1Be/p2NGoT9YSecYXl+6H8M9E9tzMYzC1sPWLmLhladMfXxmm9hTJQyla
cxjbpUYpn1wIeKXgtAWBMQN31cUx9WBDf8yecnoeH8IFxSESVn0WSggYwH/ZJV4zJpzEjaIUwHAu
SKTXjrszRciG4NrrYm6+l22nCk6Cpyl16Rp3V4PQmo35t6xt8FGx/Y3rpcEGtee6SiA0YBxAETs+
vBTVnEU0fzdct3BEN0xz3PFH+I82ulmOpnOe2QRX7mSQgSn7TVZh/ljuysrvgcQH6h1WPQs7JoZ/
QLGTcRfnrNrYun6aF8/IcZ26mPiJ7J3JwNuIylecSM4bMyuErgOpFUK7qVxHB/JbWjnX5RgITHMf
0yTREmWGuolyjkhoxWGigarphRk9GlYcfBuWYnN45Na8+WmGeLPlhKfC2mWVBLP7fSIOav2gpd9K
kHro7R4lfY4/1slhWY1vNde3M+VN87E9yTPuxlXCELSARNEHhztem5Y2wluN2CtWkazoI5v+TZfG
/F/Zi6ehuDnttE7AsftVNNupYrnwSR+hoQ8FP8QfqAQXJy9jAp0FAMDPP3Yjpo9wZjXuikF5AbfI
/aBQS9XAY5elXEiD+TznoY86jjAXXF0bfKM9+KmH7tqkiPmGgl0+Z+5DtS4CydGZpqW5ca6FqSDl
7PfSqgL/JvCV64aHHFlc+1j0f6bC/3HIKUPxSm+QuAxWYsBMOluegCMQH5nLSUOVM5gQH5u4purw
iS/ppgIfn19N0CbZWjJ9+rhkciiHKn+8tHrXNX3tv0ORB0/NhyMoj+VqSMXnsudmvhRfI5yCM+AH
yP3AQksm4u+7D4cpkpTreG2c3MntAEGi3zw7W7+dd0rPsVsIuPR5FRXe0Khxwkw8bFIXYkC54+V5
eGWevgtCqYPquU3Vx7rrV3O5jg49uk9Lt7h1n0OHWVAHVvx1WqU/abClqM98t05sxgIYyeVQIHPb
4tYinYynsIs7vDrfIwPehm02+/hEmmz9pR0QDb9vkXgupY1uACP+TNs482LryuvSeRsM+wDaqpsN
niRcUrBkVqmmrAsFnN4Mv210M5nDR6PPqL4ZcLU4db/gTTFAcQDUC6b0aJKOQaTNvINdGzxCKMR8
mokhP6AbGXcMEFjosk7BBmz3M3owkHblCSuxZWsItm2vXmGJLFmUbrXWkWERJnWa9z2QdR0iUL1u
sVo32SWIn/sQTwLKpNovZxyLOL8y3RRMP5FdxPGOQKKe50YbDK2A6ubkt3L9GjDSH/0MX3DpyK+z
nvAXzxS0hLqrKKwn2e3aLGiB2LJU2Uz+T7F0iIvGqVJmqQ08zmGOFTXDalnj1/C6ZqlL9q1tPrhR
/Rz8NP/eE4gyS2qz7qpuXDVftFpdRDXkDob7b+E22i0FBWcmch7BCJpNbzWCOblfqf1yTRC+qVsM
i44J7Pn+Le1xJJoF/Ssw74BLvdX/EIcRTgTsb/sFt8ko3bFyxXOV36HvjPb1HznrhfZ1C4TywI+s
Bs27agmKe5QekRIaZ7Xqo09MP3rJ91uG35Xgo3mw6FAKYGuI/oAXeBGcEAbfOE2bYtZuh90BXjoJ
nwViUPsvAW8rBhhZmB4qQ9lp3bec967Ab3McDcyyl0nIoJULpoFWRdbZ6cPhpOrHP9A1CfvBKnHR
wmzdBr5MUL9fRv/GMT5WUhhHSGRBswH+Xy/N0P+ERe/M7IjHbSJT8NPfTEo3n2PXJfygogQGZn1/
O95mNhsks9P6jExJc48hPNdDLytx1RclqsY9Ja4wzj6tF4Utdj3Y/tzT2Hj2y9/MLulZkMCoIInX
9tz7WKZ9zIESohRUoxeEIkG3zpPRN4gsNERz9yr63Aw1elOsv5M7b0Df8p8byBsv4pgYswOKVCxZ
GAoVfrMCYdJNTOPICafi7XsTbNnPbO5p0fm02oGh5ZLSh1mMhpZW8ZrjRNbGGVl9jfqHsrU1Qdr2
XYnqpJcuZBdCc5p5rm9PstDdkk64mKQBKIE7/zoUtO4nqY3XNKpjwdshva2gVymkB/koKJ4cVCtG
/9E1vrEg+/3C3jz08RViu1AVS8NfjwHjz3X2Ky+KYR0o/x+W2CFmYuRHdd7lBuaVCjT9uGRxnhBm
WDB9/4FK7ILwfe7cwcV2HZYaEtKYpT6Da6jyY27vvAykVEORp4XbJANo873IOb7cs/BJvO2Ytp3B
vs2oHpu/wJJoRGzMW26KcpS/hpyRuvifI2e0quW/z5odl7pn+tGT1K/Hg1pyFbbJdeSUnWGFwcZY
LR1qG/aueCWAlPpHtJebyQmtmCGwsN2I2f1f4/ZfXeQBhkwEz85gEOlDTtpn32xGIWhOiRsj0cs4
gafdCC2GFT40OFAAuMQHl1+YDtYc0MpmiSKQygiAMaq0zN+d8/ptzf0mEpJeFGS8MK96LotMvN2B
eKm4l6ZXgoefW6gh3I/kugRdu0iORzMNvIBnEBb03NvZKVf0uhrEeP7ahi3O21cjQ3aFQdLvMXMd
7bbrDpSUxX3j0mKiTwr9vXkeowKiWTODHzoMacsgOlwfFkQHnaznAsveQa/jAkzkymPMY33h9dYi
yiNZu3DmhL6q4g+prKdO083bkPPdnB7dpDWsgDLHg8XLiDNDDWp28DQ8vKaF+JIQz/ZwZIgC+PNF
FDYfaTlmHU2JsLAv8ngZPZP1rluOygL0ymq3uTPqlOGBYsfJJmuMvUo8NUP0++btQFUJAkIKbNlf
TVW6Q0C8FRwAkr6wm6hJqS43fP1LStnDCGqU9lFbUOxXTk058PxV7rCUIkXoxcnue01hMbvqHE4T
b4y6ySLjTJ8uLSihFaVh2EKCZy5qmIg9qWM5PMyF018IbugwHE9t0J0V9KL0QUxDK7txahn3eeNk
+i+l1zFx0ksvFyL/klAaFsADiMXMTs5/ArZJbcV3n2sdexJ/LsjYmfbU6sAvw1/YFpVcujtVLgET
yd/ANb8dyscZf098Vym8hWCAOkl9z+a3xibuTRcJUzGyB4LXlji6odrU79+zxW9I63vK1fTSqWUz
sfcQNkz2iwTY3Uc9kCR2GPiCMPIp2GvWA0phOFjSEEeJCzmcvhN30TTgt0fzf1NppdRMvqSV8pu4
Wjy6ObmlYvYSVTZ34hv+zhAEfgmOFq7BeNfj9MCKLwpcwlP1g1q1rIywzVQQxf63WOa3jAI8TDAv
67hVX2SeGjyz3UINC+51LR2rKBd8ANbK6FtDl2hbj/A5tA195JcThNCharb34+910fjRaF7uh41o
+eQX5BOITQJb57Q5TUx8r02hiP5h1QhIIlkYRnNJOwlHE2UhYmizFYxyL/pnBTQG7HXjqXrB+IZ1
k1xW1u8wYyNAi6o1s64xvz/rYejGGm45BGHPtHRYLx+/UEHjraUkQUEaP9F9FJyOzsCAIpIBYOQd
5P8M/SK45AwSXV7PGkkFpwYge64o2phg6es1DWHJJjL131m8VNpnzJF4u04dswBCGqWSpw5LxLW6
Y3fzmQDF8/iwKSum/gRxLe8yf3ea3JImLWC9EqLyztTTP3rgVvMTfhk3HF59eM1Qw1ScU8tmTLJv
F/H4zKdRkj9fboY3tb1nLyaNtPEhUKcmasRXxMi//md7S9mrGnxANsIb6Bjx38FgyxKY/7CXPlgE
+PI70GzGPaVRi6EUM6fK1CzaibySBvOPAh4bK8sLbW87w2d6jRImtu/gqMdrP56MbKAKicxixRmd
AtVxLKUlsS+oFEx5F1Pftp068Thu+uYE9DAIQ82Q+FzsG8Mqt6+vEEDhvt2YCQHV9fASeDZQIR7L
H478VN4OKe3v5IBXjyPGRA+0KkIeQkIoL8+N6SYpxQmSbpgn9Xe3dDtYwhIuCKoN4/POafWJ6j2f
jLkOECw5IP8E5tB/0SaWC6iGKWFmcfM1Q1NEUuONL/xjpp1YKeHsUElUOLP4RPZdDssQv6/B3YEn
syX2oXNPuZqM971BJnxkKZhw2+Ub20GZDsmBlu4pnOo8HlJfTJZBykPE8ITEapYJrD9DZxPfNSRz
k/9tbjUIbo0XGfnY9xUGaA2lveuTPiS4YZ0ODDRGKmmVMISJqn96auvpWRXmsSomD0zGFO6pp9Mp
l1AfIrZH8gmmdl8CQCNF+pb9oGKD5Ll/fFubA8cw9Xf+cTIsbRbCQw16J+EUsfu90fT6xpbDLI2n
WokL+veybXI32PxW1nx4Jlg+apKDm1rkE2TlzOJQaT6h04s0rVgeMaTSY/w4DFXn8ZZhEEhG7guE
Hh2tTNfDQQTF4BWEoWHKuUDmt+Jg4Y6E9Ft1O7nXVBCik70sESEiQBtHxyVweDUGhU9JrwUAArAo
YPKif4mSdLmrGptcLucVCIjJQFJYEidv9KFMa/Ae3OwPaIoXckpbcJ6TbpGg5LRPxWcRtfRpnde3
roODDe4LFRmlRvfizvrmt5J15dyAjiaoJU/e/IScquBUhvN+RZ6xVtEz921VQBLIhM3jwBBsE5mF
DHc39IarvQwdL5TGaN3z3Iz1MKPuBSsfHFT2YP/Mt3Ex+ZPE0yPXF7r3Xqqb88RQ6aGImNiJQXDY
uyqB7Usia33lOFFpof8cnciyPmX2ZalbHe78G9IkETPz0YhfQJislD2lEl6cy2nzIwWKbSV/K0mC
BpqdVOfCOJOZDillRavq2528sdCy9Ns/yifJlaNQYMpQOklDTQPGWyb6LlDdjUlUhcxV2O456JfY
F9fLr7VZUY2Klfnp33G31PzfqgYny0kxe3eFz4S5XoiswNJsytC93ONbIdDTscnDwA/YbBet12yc
aleMhgEUYdgLY8F2eH3aOnrwQfhbYFn+o0u+CtqsyeDRpNvIghHwn4yfrMKYV7QAFlBlGOQlC0YA
ecCkxny2s4LOCI6gGN99ny3JmbLFGfhGHJuGXlVrp5eaFeXOsjfY3q/ATUkGg1lqsuN5tPoFVk4w
//wonVmvCn6bkjWRYKySDMx2ZnC1Y4KDFmRkqdwJA5H6dfwqKS0hXvia4E3H2behLkPXBIgwCc73
+J7BKr5xwGHkwaqkwkMnEOLApRu34+WT/h9dvUSaubh+gHDPNa839pnKByOOlzXRATMmhljxnsnV
cN7xxxLOTkUMc/puBTwg7AoLc5mPZbShtWCHd4VpleL8KKzxL3smugmi9EVxUfOic9IRO2PQWQnJ
wXsrTI91PAnHrd1K1uHlwhzfrHxl+75ICaab3GB/DgMDWrG55M2/nZubmYVka4+FRzSAL9RKlBYl
c07LwTBfiJ3xoUTPkIWikctv+sVGtJk5/CgRZZcvNyYWjzZZ3i+vVYD2oyqvwl8ERvKL9J9buRWb
ApiBtWw8EdtN8Ic7/bg0RDK0g8WhoRg58NrHDCWS5zMozFKdA8g9ok0b06vmJENHsIAnNbqj1EKm
5t6zaRR165BqMrnoyYgyRW9DjOLHydXa6UO0uPZQ+fMYvPPtOjv1DB0GAKSJHDTPBOvP9ACv28Ew
jtEOoTAzLgXrw5qVvEn2hToFgqs8TGI18mJVokvhHYtlxCHEi5vMfgp/zJTDnDljjI3/U240ZxHW
xtivhRG19KCxNxnSr4af5LtriJBVxlOfYD+pLRdS4VHYUjZ5XuUa2t7Z/IaGFKFEiG2NPxSd4r29
pBveGyL6DSFr6xIZ8+vfmozGr3xx0m9lgFFpYZ8eXlgRkCgUlAM32/eDLc29qxbkQSn/F5ajGDt9
CcQeKm0QI0JafoqUlJS4+hggSkpNI7InqkXg08aCex5MZicRis6OPrtMAyS7/SGR4eW4QLVihkAw
jXBFIQPAVYbKcmu39Idt9MlwcBwJOizJ3K0w5oEZwz1+hIuR9y4kzkgqJ9sMo3bfyedfPJxz090j
hp5Kd86YaT8rbYglZcZ1lCTMh2nOmLd23znZFWEbJPoimB7QFL4JcfoBP/rNw4a8SD3xPRAKJDGV
gDveZ5S3yCCByLCO5S0umiv3zapwm5/Cladgm0Vuf6e9qbeIJ8+J8800XCq4ztVYVlUHX9tjiKc1
zywIxdFl8U2CFlTdBvQHIbEPu3RYMCUP878fQuMXSahyRAshH+7UlVPKc71drygijdVBu6Ba7XJ9
x/g+mzfTDkSyG9ZGEhkXHTXH2Dew0axxS64AwHymsOy8ZCJRStygfLUgpbAYZ8mnUiOXRBXS2BDl
kZ4KvIN5tiSSDkxZG8jpFq50CHcHDc5JbjG3Ub0X6T53pjeebcrey/36OArF+kxSQlOzO9oDQTEC
ElCLAITqUXCZGOnAx+s7yWAjaPZC6ABj33IiU09PV6H5MI3cYvAxAVHXggU/PX2BNsnV/2GmciuD
+uNQa9l4ppC7WJ+sVXyW9PcHcX1TG/xHpIHNIqX7A4D4Yhv8NTEJLfL+oAEF/2duEkmwnsrKusQy
m/Tr/G7/MD8kxrkwjliVZRa+Pncz9dgN3p5UAd/X3RSU7Yj3kkEVTX4iIuH31jzjttfdfZxCae9F
V5YU1UMIk3FRomWJUIu9ZTakhFmaSGLZnEcGeCUzIHoIlTbr6f8or3Vx5B6iKxonXH4hLNlrY6f0
xQ0JaZTy64leefSoMaExIsgSYX0oJXqjSxXMyo1zsuM5/PNrWhbKV7XYqQtDB6/tGuidxv8sXU4v
XEuhiXocei5quJASLcIPU9+QbVc5CkF7a/lPoB8HPCY44dg8USH8hTNJsfoThYz6nnCbXB9Cd80V
3ci9cYCWVO7FaYX1Cmd3Z3PmN+PXs9MdO1AEN8IE99FLhT9dDturq7AmeVlAmMRDbHkv5GHCNBml
lstCBS8nGbNgLcY76Rl8auGwuuSP79kxEPGfFUy5T5bzeav9uRsuxTJTUx3uTBKTN3C2KPTAS39I
XaNWM8ifrM1I7ryKoXf3VY1VWzW9+YJ6qaHWEbz8neWtk/+/ZDvaoAP0l5Dl1J7uAQKTn0jhp3eY
wVSLM0x6xEQ48jvNUfTTHTM2pHvD26XCIpyrmB/68LtHy5LAUyft5E4ZlDefuL+ER6bMkMHXSIft
M7nmfQBwiUZbe6gXQCXBdW6WsXxe58hTlAhid0FQM2CVn/vOvzfcZFxCeOUNVgrpPxgDGPcAVxYw
QpIogyHZ2Nu9F+cMimRX140fb0S3N49vBPIeTNwevJllJbdI2hbO1EvQoIZvHHB9gvGXvCbKApDN
mzNv/1AcCvunwew16ekOJf49qczako/xOT7L1gDrJteEjNkqwZ7jUVxwjWqXbbk5K9rnbWuihMlw
eqTuF7v5OQOn6z91J9EZzIXNyDl2vNf91yVv+ChXYXkyCX/I7WCStFUjIo/2yz894MYxep6AOEhv
sXWfflinibSrNHpDKmZ6KiiRtYn6Ydvceaub7gOL7KkbeGo7HVXakvTiOnNiEyLSNKkReTp4CaCM
1nCvnoDo1H88hxcnAQzK+rIkf+auXVs6ceDwrsP1OUJ7UQVhyTPpcCgAEr/8876RcJvXJqZx7HYK
kBmBwTWYp0Qm81M3RS1/oCrYt9nSVA/p/lLibvdn2rK5D7VOh5MdR8UVUuIHaJtkrne2x4fcn/xN
U3wnvuDMD52n8tnNoCf2UsAgjIsl0Ec+szRjAERSFBxBaBFDr8jtcBqbMTT+uGMPCfr/eM14rXbw
tuqr2KpZxjDi9g4WM9nezou2yYBK9KfNMZgs9YId2iqR3xsB816E/pvANwdNA3q1EPYID+eZ2Xgt
wcfkDp4ThsZwLv3BqgNpdRnu5iawTcYYjAsWSbGpzWa3vD8J/dzPA0rs6291UG3er3WeENmpDTsl
PbmwHa9nV85b8vLAxufTLNv8JhsTBzOzCTbiioBtbNUBhSI04gp9DHT6DsOD8Aj4O8J9YSK0hpaO
YoTPH5fDFLaS+HWXD+C9xHRzMABx1bwhdiVm7EpYVnzkQgwbzVg983AHVfkjMUU1rh6VTJlTIW+G
BWfT6fuR90uLIYuBuTNuZTd//2CzK8Q+3hfPZ+jykMMOxn8+CGqPnTvJ43FCmDkN4Ifagd+N+TZ8
LNwTde6msoyTONA3a23dlKMeigFkPSM7JpVLo+g0OcmVZZ3T7uB7lwEOwv51cHvVEgj1GyggnwSF
HIDxw9Ef4nP2Ha78dZh1tRgGvblsuV0dMCwL6TOwKxVyMvUK9HKvK5GK2AuPKOs1HRT/GYqqq1fA
FGpQRcMhr6XvX6G7gFcyjW34lRGspO3qtNdsRKwn2EycnqAdi86LnpcLdxYOYeRhLrZuAovkpY2a
0s3PbowPzpdbfNdPjov8xr2GEJZChDM7yThYVocoq6ihhgh8SuImV5k/9zGTAvjZjZFAtjxRNsM/
45nJmdk8bHA4+RokDZRuZ+zuZQxuyiVC2YZh+lMuxf7fv0doJI8gPCGB2lSie3T60ly9VBdlBTru
/B//ejSVxSVutpjYb+ii14KMRuX1GOdPiV56m3XWmM4NTGFUOYvt/pLCeNtilCljnXy+3raigeFK
u4I8NEl6hHaB1LyDO/Asd2lqlTZFNT02HwhNcOBbwtnivHZckiS6gGGgjgoX1SbYwojBrvhS4AZb
2B9VmRa436eVwMN7fXoCQ0hdeqfRq94UH97RMlN6ruzFxBXIJbdW2LpBgTMO3Tabi7Ps5570I9cM
LertlIg1jtcTHAU/DLS7iYO7eZcuVETzRdSeliEskXD+BhkCAo3gU40WpRF71QYGercZ1mmIdw2x
HCNwcFP1oymiH7BpkU75ylZGYHZNZMczB02vcLZVdM23+6knOEoS82tCk2GPbP63i7VdvkMEbBXE
Xl+OwSfSkW3aSYUzPI7buz8XhCGeJKsjwC/SMAyvMNcEMdMWH8X5t2099/Gluz/QzxdmIKTxjibr
c9JxoTO917B44vU3ExCpwqs+/mHVQb2Rrh9+gbVZeG/t9cWAU7EhDDKA/UoebnRMD9wkGv1zaCiI
mJvhK+q5ikjc9Lw6cZWSX9ZpzYSsU2x377jxIR7IjQAVyC3tpgCbAJMz6krVY+IkpT9/Fcot+7Rz
A6xJsUI49+7Sx7sksWsB11+4hhs/FoMM1c6MiWFXW5yLhcai6IrPttTwTdHEM4CRhqvBDxoFsHi+
Xp5ttHT3xCB+BwOOyi58Gb4wW4RGiz5yggCsZ0flbASIXWOZOeIroEf6H/p4p51UiIqZPFZhHc/h
bNZKJyJsRVrBz5cgTau6gN93dxX1ufpz5O9uybXThDK1MCp+SYneXZWv4x12Vd6wJ+oOmxsGjipW
fk/cAxZ9btyXRbG9f/YcZ//m6aOtvvlUEl+b2JE0HnqrG1AihJjSbRIU9OP5+hSjaHRxyJhPsWv4
/9JXh0icMebx+IXjAEAh9LcG93uH00P5K4/UX02BrAmrDBKlOC3h4hMJAhkut9Z28A4NSmdbLPbz
Jeb1KNfg6Yfe70amm3/sL5v8I8JKGnSZupBqNVmdwnQDLkSkRdzm9DTm1QudiclrJzrq2XIjwzts
T56FRT5xvfKshFyu/HDF7MnebqV0aDk5O3IKd+JKuMVGMRNc8s9sSpk88qKlc8Ly5sCUNSKVEv6V
weNif6SQLEeyY5OvJMDSnyY2O+o1ASdS1XfqHqLBu69m0vHTiQwuX7itESUvnlibmkXfrMu4Lm7R
1cRLJdj14HUc4xO+XeqDByYEQPebUcxB1X0H75T02AZLvkj4GCJEC0kbReozIgTk+h4QBy7oq1xj
XaJ8jHcfl8LfOlkdpEQuniiyFpcDxWKSTJawFHFOP7jsrTclRNMPPdpOzstnlVIaU73Jc1cndz76
JGd/h1hYQ1kZTb44AIwCHfeVd4qGzRbvfrf2XKP/I9yMEl7fLOcLKliO6wptIOIOezDzb1BtPS5r
evXpz9ZNDof2UiaysIYIyqJoIM6IHNUU7LobPWGs6St9L9heB3lBBdj1YZWvh6TNv99MojVo8YUV
FvAgIPl9m5Zh/mDy7pMCRjJVoKV1TIjvuWhGJe1MS76GmxLX7rppIgR0M6/pf9RHc2sfrD++GgBF
xLzolQUQRhHgsoPGNnS0Q/gvkgTE/RDlYMBtbSllu+XTBC0wNntcmZYvUCRsh07+g6Nax5zVxGNM
sMcSZHiGpkJsih1q5xosRY6w+PV0md/Y2ME1qXj4Qx9aJ8B9HAJKK0fHZCkko45v5H2+gNwXRh/f
4X8l8ilN6abg5p6JA8w60UgpiQl0bxPdxcahuLWO0Mh30ZDKE9nMGGpZ3/f/WnlGxadmcfuNULUW
/Vsxuwozz3W77CjIlV62c+szG/JhBx8Krr9bJrjnGQG+DgV81UT0s9gyxKnq14UFwN9A4XZrSZuZ
S5GwhInm6Ga7RJinNMYLiglh7f0cg8g441T6BfioRFNqJkiSqEQFusn3vmYjAMyxaoHeyPsGFPln
MUIlHjqSJFV+FcAkzMeGiBJzagXOqGec3zvuvtbU13Ui/rVFpLOSbPXDv7zpYfxvaLHBtoGlVYsb
f2TN6dA5KIaItNcEL15tbPPj9i68O2vwTj+XaIOCvHnKbzmqI39L3x2M+djxiLFWdeMudPw680QE
F1yBiYDraRUTSynqiiOTZAWzJaulgE2uIHuRNjEjNLBp+Xqx+C44o5eBSuPxEfLAh5Onl+q+mus2
P7P22Xxy5st6EeWTNJ/S0lxdO9e1XMqvDyKenYIlCU+9iB0XQJQmbJNhFheuYxQWFf/DMT0xQfCL
WOep6b5krQz62ZR8gMtKx20jjnV1Rb4E0XvdhNYytbcd6gz8hJpe0+69ULCbUtxC1Nt4f4/6+GzM
bGgRy/6XSEAsBlkJFzOx1dG/4ibpG3HkqjpMVlQL6bgLwAAaWNRHlt3x2RXLt73VazaiWqrFPrrj
SyDQkQ5jKPyZeiAuEsI4L/Fqag9OeEGT2B9Q2tmNpbFZy52gQJWK9Vv3vO8x/ZaB9550BciKRaLf
eHmt3P6Ufrm1K1M2pqz3y6iA6frBE/8AH/n1Mh9stXKfLohPtqss5pb8+9toGYyd7JjuvN8IUOEq
IFLtlRRodvBpzK3b3kwb7dEVKqHHc98XFT3ujPAkYslwgg2ErdB+S81lM0G7hE2MVM+elWoqRNvB
TNMh8Aoez0nDKKgM9rF4qOCFGVp5xaJmvWSVi14+NLorN6FoyE4+//hDjX+1Z/IYOjlqcV++dHoA
bsKnnPx5YH5XsX1ikhBZazPMta6zbwJYSs4QFYcw0olvFs8xER04qj+X9zAnIBMe7tILlNnhPDXg
rniSaGDRwkCEQVYcGnjIHNTNdnga7S1m6Vfn6ubxtnuNxwOVEhRNlkgVsTU1G+l/X7bHQRs2SmoE
c3EroAQ0cClJ2v3NbJf2u2X+uwsXDoD4MX9OtqK0hJ8QY0dBFDTN2OMxPNxeojURVBV17EcezN0l
PA9LXHlYHhUzAFOX3gSuA9jxklOPy6tHFBe/JQHCulD8iRXia9eRxvm9RRjcyZFenME6QE1rQnWT
OnQoCDJHwEJc9nvH4JEh0a5CegzgayfhkCXd9qDPQd12TUbcU3CLmCkrtwBUxcBfSKF5LXG0axku
EB1eQoX0vqktvUdqu2TufPAwDy2IHqRXhxvBORzxTc/jWFZrEG79DgCxU8QkdR2DzpKdksyYHxd3
lS9O8T6oe322uMmTNERHFdC5kLw7jMYa0OOFE4jckQBed1JJVQHuNWfPXEnadsH8Vpml8MbCoYgV
zhrh+JkRICRYtBS6FJqMsADfU3R0ppEt3m4NUaTGWplnb1QJEVLgP5Ty8wXClnPZuP2V1jMAeJvB
Zm+vHrzF3x8ho0NuWtxCkdhZrNcpfCXMwyQZnK28/HyGDFJ7rbSOLxI0ZxJjW8R82bJ7LOvqzU7w
3e461TQp3nmG+JmXpNzFcvexmjcOv0+ym2hrbcEUBAFjzihQGn7nVqbP0X0NCokQ00H8g0WtkR+5
TL6Oketbd8zMfF4Do1mdnQ9KZtbtWNLhMmq6fZ7aeNrbK30lk/XmAjFDTyQJoCkV8x4kVpB84H8v
Fv9FUdvgwj5uPfB2Z5xjXyh7KfbM4ZYOddnG0sGS20CGnrgtcXy3+00w8vGIns8m92s2UVitimEN
x6r3Sas5gwWYOFBlHd5pZNIEzkA4s2uLSiXj7gl6DVjOG2Magfa1Gbr6o4akJcTIQfuektU/H+ZQ
1NtUxTe+BmVZW70nEgH1AE2c4mkdoCnKId06Uz3EGrydsD8Y5Y+6HsDFpelK8J9c/i2ZSgM4gqFe
eN/gQ27ZiDo+v9VjiU3HXB/27R0KRrBRh3L6gz5N9tuUbOg8E+VpzG9Ws12WKZoB+a1YcHyW6QU2
Khqgvkic0D3PeGWbaA68Gl5Tt7YBPCJcmBBR00YVuSIq3OxhwDZpOLWkD72QwJSqrjXE9U0C5kBp
YoM8107Ey1dVPU+tPZ3+pwaQCvAA93Y64OjoBzM0bQ4NpN4DAeFd1iKyLXfJMQUMutEK3kdYwYs5
xgL5lbS2/1tZy6Mo7WjMdgZjbOws2uu98R+XQlNxl9i0xMh8PybkMOy3br62dE0SIC3tl+UoTov0
+G64zhExsnW6QGmAV+LKBKxVWi11rlK0uisMGW55Dc09bIYm3Y5yjIbtJlDFqrvXc4HNECmodOTJ
Pr0AVobmxP5RoLFxzQ2g+wlUb5LCK8iokbjjzYDQrSTtJDqDkKZPex0jjABBbU/KqMTlZkz76ZV1
CEndUm5fv+s3XkIP5Eu3Izmyc5rGJjLWF9OKayKoTDYEIUWKEAcO9H+euwMEX9P7BmUmg6BIoXGL
ojqYD874gPKqHk2g52LVplhXLnD0915ZzQl8CdI1Zk7ILi1Cn7NZvCiE79TIUDMC4MqLYXy33GVB
thANYVRbT1YBrWFzJFyLkQWF/r59PXzhmYHL64EF8e8ayvj8q3SyFnMh0PmkB4eQURSBgXqX6Z3X
DS9/F7eR/qdpSmjPXKQ2kbtkccxiYvCHUcrx1OBMatYdtc8a9iY4fVSCP3tg2oOjJrdzAnu2NK0r
PWoxU+LFqi4dvRDB3irTOmJbLlIDi57RmJhnN5LPXqdaDwhDLg+eefnIl0oAeQCayy6GxqWJZV2N
Xemir+TDP/PLKTP8m/Vc+5rxlggjqMN/+UusP3yldLXBVoi5YUF3H+eFri2Pl+E9B7uUK1VlStPi
3BbME+z7KZUobPf26YueyjHJdlXp7ivSl/dWDP/LmbkT9+6nB1glL4gYQJt1gBxr12NR8VUNOnkB
Il77VJ7u0duMcMVnG/6GfVIhl/Tlg1eagw5Mfz9zuRK+rnPDCCG9Rb/YN8ElhKQZyDmYxblRARGN
jIMWA0AnhwNaE4jrtwmI8yWYZ/Lte6ThIRMGBkUcYyySIEajQQmx5O2XdEaET+WSzfxwzSUvMC63
p2VaQY/67Iuj9HDZ/VvYKVL/AhjmGV6XOhGYvorfpUg1FiJJO0wijjw31lxh4inYPcVvqNZ7sO2z
pFuDtyaUVM5ImxEQ3WENEH+872buCavJ9i80t5aM/YyBvv8EaRfnD5E8oTExLlGsDY9xnegP0YSt
NeZ2pPuptfhEnyUIalLZZL8aRqKjOBjFcwHsz3PqPys77DnYN+boZu1ld3Bshxmn3ZrExUyx75TP
ZUp+TPaoKXuV11OBCYK3BDqBfFuE+gn1QrlaC7g01ll+P+bNFwFkJ9Hof4ptf+k7LEoliN9fKqFx
YX/BE/0PvprF7eBjCx3uPZQT8icerS1ej3npjrvbPFxakgK8lomLa7YPQBiRGOE6zEtG5mRJ/0io
GcoVgpuXY1TR4sMeZfNjCpMlRL7j3rhPaZoTHcuYMntuZaolPYE27ORes9kdFkKB7ptvVxPxh9Qd
/VGfV55YX7vUdnt65wNWIelHCKJAsOd/OcSsaFKxnfB6IWhfDJpvP9byW18UcZ0Qyu1E9eTp0WDB
X1ONQP0djk09iEeUbVfJqwQ1g2xZkGi3vJtMMWty8S+KACn5GrSyw3FOmG/mTIvPNKUfejgpCUNR
AjA0b3VqOvIjLHlwdE+rPtWe3+sExUD0X7hHbH8sbXndFvU3M3IYKrK8WdWbkwvGHGoTZ1BNG3n+
kfjr2p6bcTEKhhO2YkeVtPpDrg4DCjZdY9NUepVlYmLETjCSJKmfQmEV1lueDA0qi62v0OvjWY9+
mG7rDRhDGTFSWJbHu0LXT3mvlmH475EpSltBZ2K5Sx3qPK6nWLm9736P/hc2NeNOTBscrbOlYjV9
Hwd1gYPhrtmTKRlBeQNfiHwnS5yTt6MiRhwNC7MW5+nmiXt61mRjDcJDwR2ZqIZqT5xbXMzYwsOv
D1oGCO5PC6CoYMd7lWyXJRCbwqjSMfa7uBO12bHPbB7WEb9AQ/DN6XfsADqq4q2tpq8AABpojWzf
ufZD/l/1wlf7cWwHQC0Nwh8b3aZM2iIp1/QOXZfj0yZAV+TxyUnEzknq5Gce5vog7WmTa5qRxbfv
HBsq5Tq9wVDMrTGO5i38n64VughD6uYqu/E9G3F6HrxTZZ7Y8zYvoPzDAqzLNudM4N+odic16Uiz
frArDH+RPpOQzOUE2XgKIrtNyneFC2d+gV/eg2WOpVgy8V2xKGNeG0wbgiM/inNBTw+LH0o7K1k+
NRDfduDN+klumO2eAYFl01LDEuAJMSf4Gfesd12BAK7qcyrq2xrLLuuAw1BDa6WyFj4TzkRUBe2n
8gyOFmd+iRvEZrPWcg+CPto/BGf1nrXmExlpuGxiIR06amQZqaU2LOn/0FEztCGRB2TOiz7xxaQY
KbyZqWrCM521B31j/y3vnDfkwz0Xff5piaeJfUhjQ67eJpRiRmqHb9qUB0xUvd+U+AXY8o8FrcJ6
uSH7oUCfbCD22xQRBPbU54Dj74AOQckxhRTc2kpJdaS+eA69yNEyqedDKC1Vgszd8Dg/xTvfPOnQ
/ttGFhPadwJ+IGCm63hFK/3roi0jSPJuHMkwiAYtS4a0+oFA/pQ8W+h1J34JpA9yUEhtJmYiStNi
ef+py4ergOgJVblfXP6gB9Y2e6fX/WzoBCa2s+ug4WPt6WkJOo1qHvs5c9iQMSDDSdMqHS5PjP7E
oFNZ7gGyfy++21AD0rVXmD3tLFKipS67OHHduFtFecnxxVB9MlyNl/SLIfZBfEGH5OL3CEfV78vp
EAUa9n0gk0Yf85q0rAAXlum3qhT2Ee9oLB72QmzmyYVFH6Q0cx17WZ5noSxl1XXO13jheYFavKlJ
ggEsOaT4P7yTuERDxLIYYczytmD5l7QjDKIps6JSchLLf1DU2+M3dRMY+Ty6mqZv0DfM9iPjwwjw
B83suxcAwr6yGEjaszFxNCliDcQGcOCGvz55U+UhdCG1iOziNsiq8lEwzsliYaAovap/zVZamsM+
1q7TDFBKbd4kdmeVDmg2/9nSBfaDhWjzurCsw4LsjoMONS7wfcGvaLzLrSx3Ml08tyVP2/cXQGEd
NNGpyu/zlB2XS3XLRPPRqGhqpPdVq537+ztC3fICPEBgKXtUYrulAIJksAxdC7cTWTRmLfnGTFVh
3iDDviwd8r2oqWgLYUT/+iseI6qSgIJrWrCP3MedrV+7jfo5cAHL8qrIwojMXiXmyvjnGkoNwCnG
di1dyYqxZSAGM1ekckFsEIzMZU0luwJb/FyRykgfoojNWpt+mEeGN0IKahnOjNndDzSAi/0WIj2F
A6zDXkbuuPWDul7pBU5O64EGzlYiZY3qS5EL3eSaBKflbTIk+KA+uqWzRpDXn/u/X2FAyQK4bqcE
PBZoTxmyD2B1cCzOWaFuCP+IND2xJxQ73UlHVytCpM2uPe+u8d+VKIN2+atGsIOcj806KI+gE+BS
DHxkbeUK3eDU4FuhWPwj6mphmDiSqZ85bA+OBKfksHAi1IAOBLSxyKIJa5WhQkECO5OLG1AHLsLW
AvHVAtN/r7f6D8v/sqrYdD9/0sps1uRkndZ8cX9LcEja0L/l0NIBhhp7mMqf/g/ftnzWF2yOacDh
N4ptTbNjE4dHFrkG5GyT4v1p1z+DwkAHFOCy6ZqktjuR14Z9ZU/4uDqBogO2UAwPx49io5vpeaiZ
Qmpne0G56h+aTdjCqRqdsVR/q64SHnp+z7WZVvlrbCkGAqpwXIBW7T1C1A/gFhq/I4RRrFUIZXVa
shdquJJnQICSOmk3d/pBRhoZVZmsoFkzEAnyeNTkf3CGedocovmgPd932LiNaoE98ksH44Vx57rK
bMK/NntMe/HS88ocgTGttx2dvPIDziWqoBvZxm4ZzBceUlgHf84TiRhtY4+JUnN+I+aAlUJjJCn9
jZMhuOUgHoi4Mv8D0IAiSmbW+6/9KSLeEjcwLYyPD9mbBhK8PPU8Rtdmojz6fC3Z+/qbxVwIq0Ve
n3UsGObqNIEjMSWiHNOKhdMK+C3VAs55GNa5VBP/Itj54m9Cpp65Tfd3cd0jKo/GwJ6sKuxbX2ut
cjLD51IlzbqTOHy4tUic1FnqBf2D27fAc38/qdKP3yPy9JzulSbIGq01kKNO7sX/zZX3L/MSFosR
GRCt6wo9tWgxjgi1j+WmPcY4F/XTlHYh2JyMbnm+Ail3+HXs76AdThZgJoPeFsLiKAPo5U/LYOFi
1ZOC7cKT1h7DS9FeqA/h7chbo+ajV6yEQOwt+tFQTQYhDJmszvmBicmMgE5GbodtvEX/lWX40Fgj
UYXhAndlOmz7NDWLfIFZDGW2g2dekJ0cbM4leIM3hbpKaqWkKi+BEFPoycrVyLjzn+r2GNc//a4V
H1/VwrDvaTVfqwuee6U+laBaKKVz4i1t78TCtNygg5azO36IQMtsA/3VfCm+I6dxIm/y34QgbJDN
SP9fo/eZ/pIcCzZRbTeWzDnrHBjbrx7A+aWX4ZvQPkEQR28BlMI2PqirFWJnBS8ppypSst7cN44p
WAe1ugrBOt8+zqyHRlF9ohtaR9GtFRE2pEEuZswOrLE89A9s80ZjMG/6zRYI52Enpl/8B7msARSq
DuElQ/BHJ/UJTGUFXtKL9WPd2EvK1ScirDxE85ob8Vy1TSh2xVTViGe3sLDmgua0sIy/jw3HlRH5
nBLox8jj8zqb1CGsLhm2Kb8jvtytgk+uvoQWSmLo3SAPAs+RKbHWjww+r4/dNa349lGsHTR/2yUz
H4a/AUZlMCexLRgC8xJ2BZvUVbGGxlpRk7HrN2stGsnvk3BhNUMFY+3t3aOarwDJ9oyKAnNsYhEm
kjI0xC8QeuOg6E2aPDcrYAtuwjpFDQmt4U8ab4W86awdz7bR/y2IW09ofTEOH3MjdHAkp9duwESD
qiuODnHlB0pYDhb4ULI/Qw7A/hDzcHZiZlcxTvM1pyoksW62iM/Ng8bIo18vGxkc7MM8t2Qnqmfj
lt364LmzJUwhUEz91F7TxzO2V6FQkl1L/q8veZ5xDbB0WZPSn+DoogufU2GKWXqydq5fW3yqJg8z
M7Kk8HS5KrFMu4xg/PiIR3nzreLi8Je6cDXjTe/sPdM8NcVpXM+SHYmn6eOdLfpZaEugFpU+HcAn
b4/ViV654r6oGsW52OZO6GLRd+pEhg1Uf554GWDHYq9CUl6VnMpEIA7Ndn9KxxsMyexCxMPZOFcr
eTESiCL9IE/yO50nyTMA5HhaOg2EdM4HFt+mh1fS8Z2UbNX0LwTWMhweXhkR/cHhwxU+2NSbMyrV
YkMBwkWUsireUPfnE7vfokEa9ohzOHsbS2v47m7cbSM3ozDAx0iBTOgJVju05WgKcajhWXHt0KTW
EyvZ29Dg6GAMNT2FMUTLvjAN8gCURCNudWstvJm1vyFPAjGhzuphHWHy1uy+oKPSMCvZbFaQEqJa
3vArfXQaoZoatszRujUE4zZ63wu5knN6gg01zZfUvXx2MlcLolvjuJVfIh5oUUmv8q1T4dd92OP4
a1rHQBKfp+WVuddxF+4FwOX3f6h6U+HHAY2StEUW5JEojEkqUQPNWjCf1iP4iW5qX+g8JJitVA35
sCHD7sWpDMhvMHa+K+D1VhrAJjvVeZmxyqe69tMcHapX9vx8EFW6BT52/m6TpNOlXVR5bZIsjYkf
3c9e18XtMvFV4VCH2PAdXZbJnjmiWKhdlDns+4vmBin/BzvgWxjdRW5Y+7iuMyTeL7zrTt07orN7
+RIJMyH3ZTkPAfczeUWfDI1r6BrGr5EedGLA/04RsOe4FcwEjfGgCJo3BGOiFNITsbojp8gc7YSn
x7hOLpmjZN2nFiz6Sz7GuWpIfCjH7kTzIwT5zWIZ8MSkpuUMcqfNeJBW1dif5sNCFnPSe4/b1vHP
badho/hNX+IK9BDBFXVhup7IIVwhP3UA/j7k+D+D+vDZmk0FpDLnNLpFY2gIqs/Jg++4JFP78KNo
bQTuEdlrEqSpZON2NIG3044WuISxFMEnKcz06WPllg+Og0RNYJoxBIXWxdpUyr4zI/j6yDxzzGfe
MdsC/VjqMzRhLntxkov4j6CR0GwYcuLp1J0Ok2RtXl8E5OqjxewOewpdpHj5jQ2UlrK7MYOHGb1z
6J2+u73LMTE3OJb7D/j+hJQtLCF6QlXRmLVroWGDu5lJxFitixJrTPm2wAP1Y+kagM/nh4CzotWX
hMdtBY4D7Mz5RTIMGA9D3ciJG1653qOQQDGYcyh3Oq6ROrsXkzKmE9smH5hX+lDgkgwlw1sEv+0b
MXCm0LscjChslMwrBqPuzEeyB81cKP9ExWSmnW3p5QcNF2sx0VKyo/7Z1HtvNeiqdViXa7VPXt3I
r6zEd/SXOVZFAP5UBYSG/ZuUqRm135lJLeBQpdIwfvXumBdmPifI/gA6aL68RTmFW0pSrEZZRtk3
1uu9mdhSS0iYAYZTtzk5aEtAPCKm8PyTqD2s5KKvBu8HgWuCZhhgiNu7EIfRndSW3NGIB+Ppu5B5
K+ZQrob085c3ack3JNEc9s3FdELz+wNfJruKqw/4NWQomLgLCi+4DytQsCif5z1PU5RSmtVgkL3r
nJoxX7wpFSnVLmpsJWict2JtoPvcdEfRY13lcnyogTonGz/NaN1dscxWOrTkDaiGtyE/gz2zZFBm
tvTZkuKsaqKR60FBJBy6+yzLBrskwLgFoic4cS8YKnw23yRU4GeULAR7EaZQe8UA4cUUcKasaqmO
+I3Jzcb7U5sETka8yCeD6L6cDfK4MCfA+slHf78qhwbfsQuvPcTrC/ffry7s62ExQ9+tGHOpUkPC
eK11WIg2xFW+eboeXaV/J4GkFBho0viEjtqkHczeGDm3nt/jcnbgaz6Qid72fF0ditOKsSFj/i87
aPOCSK0PzaVD2V4ah7kH4RTGWcyuNdxV3Y/M9BDgmoT2tL+vStEhw1GkMbUyBVCXq6vYygSjj7QQ
UVkoGbnFAlerfqDahG5jGCLPhi4qKUeNbUnHPuhrs40ks0glWHmK43/VTmCpG/YvWq892yb+lMjX
qQGbtgmTzSQl+DtwT9G0s93WfAC6zFkKN4n9T819jyJCJyPCULCD3H68QHxNzORHT/n1KAcfuyhO
sy+C91AkLhytCMhr16A4qPM08i1MTxxC2HEhR/bhP8Pg9h1AfTlCzeHqpyyZ5/X9Dn1mCnbjg17i
Nkjmum3um/+L1tGDDcvvzvz/+OtpFBss2Qpxd+pi3wS9moYawe57LVeMU7NrYP+v5LE4MIVp9IgG
CYtBZ/um8JEGoUdoUCkZF7X1BZpqPzH/pot5vLK5SxlXnJdfCfBxpD6rfb+QJRtrB/HfpgmZrJRf
bALq9eBEhA3pGy6tCur9KQqQ2DKNhY/7GfV//iCNyqqSYEglDhaKkfzaGiNjt+OpPmWHXCWWzNph
vRxFIboUBYlgf+dKyC7vdMv9tHXtjhmTwJvTr20PFp/0PVz8HvHeTdyq5P/xbBR697viNc3XAnOJ
L2LBbr1GEiWwJYbgNmf4/xIfuTDfxjgBV1QWO45NO7a0JpjpZkiQoQD3HjUmo5g2Ji6PdiB3x3ke
+rAvDwjM7fLl1M1dI2j4YN8qtNbqD6oYn5z4H7OjQwKR7J8wFRP37ghc4dH7+G32Cpj9p2zeJoHe
sbwWg7tsc35NnjUEGAp+4lFfQQYCMm6+4lUjodoCxTP7SDucLPmx7gVnbPwAMPlVLEvTcc6UQLzk
WBo9d/NFV/qmk+jUDfA1cpIXVx/+1kvNK6KMrvYeuYjNUVaQ5ZL61YAYwkzojVTnMCLPLLne1v83
wmv8ziPLp6oqM+AJVGQibafS03XD8C3OLlbDSvnZxlE68QC2xKwJSmS5UbmBpiyZZd7qEgoQWARU
7ruo+ohI5+pP1qb4ZU4GpGS/DzP5Ao8MBiyjRHP/6eZSJg/U30YDVtNEARI/8uk1wP0X0EtJ+Jps
kTqga09P+d4TzBFnSD4WdmSEoBmFsmiu2B/o3L1wbYCgCrctpShQ1N1657Es/aRcaR51+Yq+tqF5
oKGiTB4DpF7xF20tam0uZWwYxpB7FCfnfwPy6DXo4Cxi2VU4mwaQg9OIa3+jELF5eInQ3JsD1aYP
P62FLTgfhiJAHpQQnMVBuZEB2Odgsa9y3htycX5lWi32M8laqGTf72SFu9StZAjZJ2wwbIrxor20
KvkcYGsTpm9+edc0eU0tiY1/9Y94ZnznIcwMtFAhPbwhb85EV+HjezZBjwaLd8V66oFh0OKifPY9
7rSgGczpVNykzwnQPkr4VWp4VtqF16AqrMXtrSPZ6k19nQKaVbxykKdCxf8ofU0YZ3Slol/q+3s5
DSBfKzFD1a2uzpFYwbzykC2D9lMq32wJE+mHAFKk7+Ka7Rs7IOBdJB90QNeMEDFP7DU64H/v+bhD
ptmqPWQu+N1hZUqlAZo6WCl82xPJ2wNFOLazfrlzYzwuAtVpQZB7T1uoSlw7dX5ioCG5x9kjuUxy
eIlvxxpEQc9r4ylXYehg6BVcVfG8qFIxu9hJ473EI6Y01eTQ1v+/FFt94a6RNhBGacstVcZBh9yP
DvB8CMrF60LwMqKtBHLmPY8blX+owP4uCUWTXtzVg+8VPaG5DgssEr9k/VbUPW371PCldK8xWCM4
LRHp6H8JFdAqeA6gJ1GCAetpQIgiCCg1Z+wLx/na2BObOaUwIGdrRlYUMbnIsFa0/u/GhTfhJZzQ
AIgFHxQJazQj3w+1G7c0VgekeKsL353H7UwQ0zJiHPta3SkzWlphhUtA5n5zlxA2UgkNzQKKKQjo
ncWNiCfWUZTjoxAyiciCJMY+oYOVlAiKrG7uFtFlAhiU8bxuzNLfHcLMkHxjfAY25A1dcSeW4qAE
JjGZfP7Z4LiowgJGTW4QUwL3i/rtk26GeIsi+AZs7RMdl/xtlo5ZEHIS3I2eRAoD9O5l0SXyvp7N
0aKGZK27KMkButbfWKHAdFibW9hYX6Ek7oUhFR0T0vM1UQRYlLcQuyg0zGumkXULN04aTW/prWIL
EGmSNUiYeD+hdM6vmxsVgReTnKzKHjJuUDKl6+QEhG8xH1wZFXK/xYE1ZROcyk56y0T85NdRMJ35
vD9VHlyaZhK1KzM3aKzXv9uaXq0Shv+sP/67Lav5E/Ra+ty73BfN9I23MMOyPcji0oVwxJfXYA21
VrbWmwXDeopGgctB31AmCKlTLHt2ydsPaLaPhm2kNQ6lZ8aBXd6VP+MsdBRBY3Y9yP589DaiJ+kj
9pHk/sXZ8RO/BYhVPKko0MiVoV1i+HgsnY4lvkv6pwXpX+NRrH3QI5DaX+NfoNXo3JOMNcM3+Hg+
Fxl4E4jR1274Js3mavbxHrE+O4GpFJPkDv2olLJinPbL1hulthCaFtSfBJil9dAXpFtAsSSjvkrf
Qb40cPD6H36kK0Rj/OGuJHv7F0LVnUwVxVKBCYX2ojs39qefQn/VujhzGCm2q61PJ/HMtLvUvNzy
+LlEgCotHLfOVCpVzUEFLwERu87z3S+lx1IErfjxMScxiopsqkB/on7W0ZUoEuN0ixeLCTFDXpBm
lTfX6WhGen6HrencO6yfAcxzFpraueNYPiS0xNOTp6rXR1HMbEwGmpuxWqMVWKDiYlQ6mfdm5cRo
WEi/IdFTySfd6W3e06I5ReuVR6V6/8ZgxdsR2AWYh3+HlxLylNuSa2/DywGPYC3VqQasfmaNUYMT
oZjqdAdFWbzumCdSEvgAERS8hsc3EmmQCaiCzqbjCbtLJd7dBHLfhUO7JI+wvzWM4j4plo5Nk6zg
/IXaOZ8A45YPh5W5GbfeoUmzBpwExJlZlIsqrfh08L9xKw8zFS6t0E6v8CryYsme9Rqsq3bvfLM9
msQi4dIoJU3s0jZAQG6r44gM8dfu9q44wcuG+cy6mkg6P1tRo6hooVRcsENPg56vrGEflZRsor+7
uklwGqNiI3xQ8mIeI8xY82BZJGYIGKaMqYGbfNeQSlTCU03IC49oOwCAKMICkdzQLvNDoJutPbPs
yliO7CXHzI5nLJKFCim6aKWFSv8xNDDuxmm/b1shFiljdQatBVATzeoUhLGJmstCl30yeS2PAJC8
/Phta79MkQmanHcVytYz46Ckqz0Om+UkpnhMWvdlCcY7XSg1vYHYZNLwNE5ujBdjuvq9Z5/B8f89
BgWVRk3czooiFPMOtViuMrzaDd5TmMieN5cYjZV2g3AHx76GjuvQp1d2qs/UnbuCwrDaC2Y77lo8
JnPIQxac+gXv2+8Nh3QgMZn5Wlxy0hf8BmXPWe3WAvVHesguW7x1caovXDSZwjvGtias5ZCOrHbH
zSGSF0Yj/cvta8EcHlzSXwbhXRMs7H9Ht3Ugh4ql76XdR1AuwildGGKfJr0m9vKel9wlu/P3jt+r
+6Dft3pGiZ4oeeDWLRdC6q9zAicfANnDrQGu+EEtPf6pZsDUGmWlpykB52n0s845a8Q+zO03GKO3
Uc/zRLUNCdf/Zw+6RheT+EyxsICVSzuS3cXUXxNkRzv3EYc4mnl2NGy36sqfXLXpqSj1PMVCGFk9
M2DuoVEALlzdsB62HTsTmjfSCA86GIJ6rgLiJDK66RMrERW/Vf4K1FvvoYXTADLKsyr3th/M164a
N3RuHXbMY/lrAAWkvV/Gcb1jniwKdQxA+MLoHNnqlwaIx9tqWXjetqDwR3ndq/UJnRr/b4HlakaE
b0BM3wIKOSDDIPUs/I/Qp1FEczmNOniQpSOjQGveIhR2fmhK6nDWdz0TkesLpYQzM2eLvtSM9MIT
DTa7RAwKtQZ6sMhLTJn7+XTo/v5fwf5SIJ+e0bnsdAs6SZM3HUK4I7Wko5bPivDALytAY77x0GVv
J814GsWamesaHMfQVAtkvEdRIQudf5tGFB+9C/si0OBQJgsUG/HupuU9ujkUFU8ih11lb67nUeBo
jDIxnnZwfFKGrVHhaTOwxIYUUn1JXGQ2+NFjAE3HXk8fJtTEAo7/1eeDOiVjCvlxgwmp9h+dMySb
oH63+kkOqDlmH0kNRaQlPkqRtP+w4yd9hTKMMjZj2lvo4j8LznIPmdDXisy48FJJ+8IV09mYU5H4
YMlzUsWqXT+Pja7T/MVxS/0eRazh41D5iVOzywLeMshr+0QKmDUQ9LWzWncfv9d/jIpL3fHuiQok
7dXcR/Yq9KyjUheBVqqR4WSr+ZxeuzdATsPrPgahMRj4pJsQmNemvrFkUhATaDkgdRFRjXhho1Uu
dmEPATKlbgd+zxgWaRIipCG+8F3XGhP9oIS2DB8JMyOzcvFDa2Hj3atoRBvrqOS+lHZYtJbNY/be
W+1Wmpw7LfgbvQcI4JtFZM7DyiaB/AGRIuJJc/FFetxW8OmLWaUqxNH1AGcJIlSnlXmZPd4z41Rz
6vnsM98eRHwaky3WPtiMVNMjTDlhTKVlRPAG3w8wem9kuOOQVogJ33AKkU5szJ2EVyfur5Bfp40/
VUR9uiQK/nBYgVz8+evUpDtbDRr3HEe8tTNtII0b3Y+iGRLKsSD9XeNj3w81vAJnv0yRYAgzc/Km
sMRJiYdUSa0/RO0+igdUC0cqEaquj99KSym0XwCHHu4U3m+oM2+aGlQ+Ynyum404bCZ0Yx5FiNpQ
WWOEJUVsmae3JVK8xkcsdoSQAzs6lSBBIz3Fi+kk9/wvFD3m8MrjIIsNcB8wcHI7cW1l2RL0wQSs
5qqg7c1x/Bc0Q6BpmwMT1JbCCmCbpteA23wkGqaZzUJcIuA5Z3R0FOO5Axj05vZQ2tKFMNZM0tKl
DQzTHeaKgxY8QCj0TnIj2MXQ2nTRO5wOnULnA5hdZ1Ud3KuB2IyiWEwj/sQmhgSRAu7OyumuXWh/
OqD8S0kLRUPf21+sRZ9L0SPW+Q0wpDtunYn/AoqWdExJqknZj4VvJJO4txYJYkKTK+/QjnW5k2fq
JDk9rmiTB8qGENdiY5Tp4brTGAPOoFMO9B8xAPQNmSRuMJ//e49J0cTucrs7stEVwz7l3zOrtKeY
H63xg6JVUoC7E9Hj02EZmbUMWYcdV4YNknUqjCwrrSb1G3NDSEWBDuzDBU+Jr1kJtWxRrbVH1Qhm
TDU07oMRYlxDT/QKBMyyjSr5W+bjhAF6QBXx0FC7Ia8yVzrjUQUgELOsXmeBUxukIoTmh7GUL4zr
VJRLAJajwOfonaqyCoOipEtYgS/ax13MW7S+jOUmcWt5ODnIbiSBoth6Cs+RcdwZAPkh/ogsDJwG
5UO0/0rOB4VVCxbseAQ0EypNtv2Y6Mdc79MJ9CiSgA8pDvo4q+w3oN/7Cuu2mAa1eb7WDDPQmQsF
nboJMQEa+eXXEM+ZJx53JhsRuCA71/MWEPX/fEVGz1mgJhto1FzjXZYhaJ5ZDiw35yAy1IAIPUB+
1DmQPYJYHfzXbQv9CgK5K+RIY61tk8xElPXCcsrtDJb6nTPeSE7+XVNxCV2pbn2ISa/oIrLY4SO5
Mdnm2C3lM+HJzzsPfJX/7fgaKPtb7tJK6/0KGgO/h5JkAiOAFQgz9U20b+oUw/BDFiD+FflSAz76
+Qr0BiKYs+CwK9TONLdd15h99TwmOQbaw9ujgdeD70DCorV2J+ia5umlLFfMgMfmNY2MZIJnA4EW
3uLqvLtdxgbtnTQXz7dFr2i96T8FEAAWyaBnfe3Q3dPiNGdYkjaKWFpMCspmOhLNgkN+wEm3UH4Q
myatSrS823sOwLgnRXQUyxUiWbFOv+lHNvcpbGHw0UW/yDkl2/LVaLXrSQvvtamk69kqMMU+C8xj
wI+JoRow/W9qMBG3gn6BtFtnkyzKFNQZJDXhy9YiCkb2qsVas8m8Qml+wtx24QuazHrhv8h/JLem
GXeySygO8gC8ykkJUWyj7Lu5xMQ5fk5xiiymNIWccNs2z83HIdKaMeK7B7PHJHPIOAz5RC8WJmnv
vUpl6pGK6q6CmVW0EvgjnYZddx0UxBRJRXvNDh0ysefci6JKA6DeiqAPeZ0WaTVaV2pPD+uJUM0C
jlBmFsssB84eTXfpf29ZCsPpw3NTUc2QulUijU/RtSRD0gH+3oZUpE8QJKHfQRKLPrEzokhQtXkq
flrs6PmB68O3h1VjBKDZ7vbb7scG0nO++oc78R96DV44CdCplSN6K/43Hx1apkmetiFyuCI3MwCu
7pegkr0bLYqO43kCXlIjHOIF46D48LQQ3Vr2K/yDW8cyxgV4dJFlpWrPgSWWkU/kYo+t30VIoYt4
Ek31V02AqnnJy9l+eU84bf/jlIYsifd8D8+MS+4ILsIFMwHsh1RgFl3FYovHmAq/F5BvsBv4KIW3
CYwc4jrHatNCjJjdNhz8ju6BDBJN1X6u8y+k0jsOGKNGiiWIvHnDJxz2+8Q69sbOUmZYK1NJHQt0
MB8e6pNgRQM2O8gYsBsmowBpr2p++mkUi3BudjkemqeEydxEvbLcNnKDT5VdsdjO69mLJ65CQN/D
DcP306/CSkWgTAg5C5wvICi0S7l25BplAOWfwKRQNifcZDGbgtZcB7pY3+cwFI5FiTv3Qr0foSAu
F8tgyDhlHuGJNSa1Gd149gmOVNXYnftxZIt6jH5iUL8MN2UGYHHUknryn9ZlbkLqElbiFKdJvmvv
umjSWM1yY9m8BhutzjQ9L2sNVPT+c2XXn2LXwxZkPshOT90elxx99eGhCUujYVKXq3q6+dgg1wA4
sUyvO+PvLP6zj8ehqrbcOMsb1ZMpVggm0O2xePtnijGzLTMJLnzwj1e4aExNjYXxIa/WnWW6ui9F
4MB2251EZnKEOgddt/bfsSFOnO6p3OdBSawMVj+3esU1IeBEBs8gAezdPgGiaXtH9KrOWjCNJ9tP
Iz4lUEtMa1ke9J5kEgccLkXWlU25JTBa8aXU1+8bSMmwyvngAMFVGXkOH3lg3CckUJArxKjlf7Oi
bWsFlFX7RCNDJciw04Hq4WY0YFb5PVkNKRZNLDwP04JuQL4URXZiq5V3jH/r0YjevQuJFKRdyZUO
en809zzeIlbKqRSAOGi/QMI5XMkt9L0J/FigL/w12jnxMb0lrWC/ML/WTYzR4gITWhjBa6ySV+So
cEaF0QOVKkYBlNcQOPhAw1GkSUhAIW8mo876hmW6LC+Di/cv/O45s/VE5YATBcfRJ2TwokNzF4ar
dPfHakZTemytHsJUFj9StPnr2tF/S8qHC4knAM4CQzdpmpu7iP3s0uVqLuuTRtutO/bJ+FA4I53u
MAL51i+xOTSfQdIReddtvkJVL8ZjixL0qcKc+fgU495Xtx38/YAUJ3zMH8b0CpKDUW/X2I5eqr9K
lmqNEVIdOJg1FC8BYCUWtcN8ufBfBVxPPsyNuxrAVG/ra/5UVC/VS4XtYTXnJaHX43aF5LyWCRlA
a7OpEjYg33Hf3QUGqIhokR6BKD7g8WSSWyOiYhXAt6pg8ukmxrlI8CsXDq1bJsfj32xO4xrb58se
4mymECgE9MvxMFYqAmpMj3+1noK28SoTWF4gIeQ6t4bh/qPAszg9EXdxdFkBFG9kq9a1MVf9rLlj
aW0umeAhWScH6uC/G7txypFD2n2nZx4ld6zQEInyrvYaoAzDhp3jQSPRvfuH89wTM4EeHSm1deDq
gpzs4152tlvrYOvBw3MydZAqloJCK1vqDIrRy3pf/45rYSrWjFzOZK+ZyS5mQPR5+JBXk+n6xSoX
sFQqNI4oGgfQi0zIL7z78/Gj1dBFMBxP+wBA5Ush4h+mM1RBniT3gmAIYpkiaLVNQdzb1GqTLDfe
SI2A8Uu2MnXnh5i8ditiHpSk8GGv7SqZHokf7PrUeMs1iAR19WSPnvXaHueIHFwFcsPNHJtv1oTm
3wW26cONdqamlI7ndk7qf/IdwPT69190x6NvUAMzx6ADBZxzAuYutY9vMuWbUGSJd5/5/tqvzDul
LvTD3U0VknvxiOSz6Gp5hbzl6vue32ci/n/uLCuIwb3Px3/74Af8qaIXt+z5wW9oaneCr3cOOokH
Tq7sScPBteUj6iJTh6S2nKyHoTl/2eJHCctHPEooZhaaHN+njNySV1+zjUJDNIWPfE2r9omygWIC
fmDGpshPOjd8pMWWJOn0177hLepn0A7q9+A1RTw5MwTZtyj5VZVfnmvX0CBVfWOj305sTRSseaJc
DUknNxFyPtL7JaGLYq1QDRDbF7dISaqUPDqyoTcLw3Pezn1t7ph8Rix2OEkECdOj8DgmFSfkh07Y
fYCOxlAPXZD5Xe4pyoz5AczTTJIiTDBxfiy7Z9O8U+1if+jpnQE7p1iGALo7hbGP7GIkFTOv8ve1
b+L8pZTuczoJlaCHmeEeyU83pFd3eaOBpO6/9FHvbRPURKUpJ6ZfMr+4JwIWIIiltV/j8rNAEiog
YCavWK3X1AwApSxyu07Lo592pE/tbZXVDmI3bAxCCWk0ygbgLKynFv1OAeZ0albN5z+pVf8JyEWn
OvlzBdywoDb7ofXea3dbASGSRCz0bee/HaMOiWjjhqINq7UE7OCTWtAbZnll+Sr4gLIxwC9ADc4w
QLazkkVT1qYideFquO3F4xuKwTTazV1b07NkqrfxNYJa8FneDtVjiwuoDmLESVlkyq7E5ELnQSCv
kJAt/MNzAlW/Mk1l2E8nEayFxLX8FV4e5EfnOiyfF+IRgH9D9jDQqn3zKAoEJchefGM1G3uB7SLu
sA8c2u6CIqxz0L+o/7GVS48blaGJ1oZcZ7S1dmzCwiQowh5p773wL0H13uWshGfBYtp7PsLMG5V/
qNi7ynEXb4mQTaBc4+HVF1E+LSas8FsF+JG7pvz/JhRlTWfcYYW0z/kGZ8WVVMMipsZgnsiXB+KN
3xljIix5W1cgwi9s7YBS55TJJ5hPRUs8Nb+O3eN/bzs3Uo6bEz3t6uiC/36mUw8j8XQZR0v92bMK
DJBtiTwn1MqfR6sfeUT4BYfBW5FLYROBnxokjuZa1NtievYdNC3KIf2Kmdxn119PLX/D2i9WLDxg
U0vCeLJm2ADWTIXEUrFbIJHFvRzBlET01DS9HRZhkVBLBb/SeK4JCpVUqh1pw0lwa4MX1i1/TC5f
cNdYkGCYRQjYCmuWxr4N0QAVramOCEpPOQ0oi3XsCc1lFqbj/eBLsGcOTt0lu0PtgCtHKAxhxhdz
c09jkmlzQeYtRI3mJ9npLamMqhFd5vVjkPQiKfuvgbaBqwLeTkQWhBovk5x6UWBe+uZSRNFoE8cR
+dvONSgCfQ2GtmrG2Mz/pp1HrGJEocrXh21LBxYLBcAk4O90fyZJKdfThm9EP3WnGBm74cgJtYUQ
qnQV7oke1l2DHFZCKgJ9VawUpeopbgrl8T5VEYu/mB1XpFutg9qoRSgTa1eaZQPoFJfIwEmQDF84
i4R1c3GJ+jjfKyjcXAeSMMYsk9v18JEayaGE6usreDjETB5RfQiUWiHaFgE2h92BIIlxEOsm5k1Z
c1zwm57f/JZDvHmxV0PRtzbTqESwxdInHQQaGNZA6OK0z2CHHXrREpL6mY2AUofkdXg9mqCwp5lr
quH2IV6Zv87tElEAhf4roj6VwM54oKUpc69mOhSVR1HJecYaicRbC6fTXFrJv5YsQZzPmLbkms9V
k1RG4HYqlmTwFylpp0qBYmlZjZ3pPl2avzjxGXzzD1ez6Jas2wEvaLbkbzp68pRHYovKFZP/pLaf
BwwXsqhkWj9UcA0W85GM4i/PO16O7DhYyYa9jYmEKZu7EVgnzolZplG0E7jzFHqRcO713pGhw450
hsDdN0C+xwyqcurDWTS1FjOKmIVgZBT0W733wUV4bb9QAbLa0YyVQjiMtkj1Iu1AmgxaTd3+obQs
q7arqs8hS7S+eQRK9v0/qE4QWurkiC41hQIG/0ByXuqaj8olpNkj8nAww85ZsPguJ9a5I5eLx+19
MlkW7nAGrqOa15hqv8FV+iOEBEwTR1CPuTCmpwA50gW9xcf874WV9NzJEIFEk05SyN9yaSDWJJlX
hyOR8v5gFTu6BTgMjgyDUt5jUX8MmP9w5QOGLQGn02vlRepRqMY/rfgY7HVN/6Fo5kRV/LMsYFzt
froVpYJrhW7i4PaYWTlaL7HgUSWbOp/rknr7jhtj5m6OlambYyB+bMVQoJasNafQfSMU4RJxAu5b
sxDs4rj/dKUQN5iF7r6OksAliIrqgOiaCIy0KkOn4VSo8D8vz6A5tcd+AnqYIieugti6SpjP8/Hq
eSXSG70KmjAJ9j4g6gK0Xz0x70Rfp3orct9EP3Ywt9xyt3oy8tBor35M0YcXr08X+6jwQOVVOjHA
z1Wc7vaL9+n0N85ILNNo9maAdlAlPw86KGs+CVef0bk+1mBtA1qoMMPbMSggecTvnv3vH09qCh7C
ZOH9W1/ulIImviXJ4zP15zpmO4xPx67mLuaWvtTj3BnZm3s2Dxj1a2OPpVxBu0nQJR0baJX7xU+u
wNYlmp2BAwvp8RCsMV0DrvgWf1zEl3tVBXnFsP5MdWmU42CvQFSMmuPdAIMSCHCeaM1XOb/KVNOv
SwRsv4WxpGwY+pTRJm20mZ7DlLy7ueBQhIMuVOjvFmx+pd5WaJHcFaHPZ2Rx5d48CP3d6G9qGMxC
990/8R2tdEfIs6oLePZzvDKlXIkI58qwThHJPw8wm6+71kUFK3kcvYoS8RSauMPNEy4OyA+8shpm
KOcokvfAv2w0mc3szl2qZworCc0D6T1wAHlHwNg+p70EWQ5WlDNgA2N5LIWlmZ44mzXpAKMUE0hs
gmUYrMC6Q+hr+3+l5l9qE5BCicCwb60iH2+bDBWhbngRIPT2c9DrktVtXhd0QZ1nWTdr9XnPbCUN
tdqUpbgjGkWJf6kVRdPD0PuQYFm+caE11sNO1nxjjFxm5iNXogRxOMj7Q75qcYyVyg9JRDjdmLa9
SJ2rWrCAYdHMj1InajHuIqT53W6hy4bmFj8jtfgCwezgAQXkB1HzvfCbhPT+LdVY7maGWweI8uLh
UGjoGctRHRh5qLjuhryZNF3ZXiIJwtv+gxK4Vv7WIWwiGAYz6ZXpfBAt3Lo27NT5XT4WkmXvTtx2
ykLgnL7wc5eOiWSBtIfYW/0qQcATl0LUXgFZoym+HRXom6zQembQYG+JARzjBiH6LMpMC89QMuex
StFTmHUlMDsc28sl0s7XcuoBCmVCKxE4apE+1BHYcdT4AJHjBmVWbUpyKLy2vIunuE7+vAObe7Zc
T+Sf8vSIQLwmprYScpS424fzqjv5AV+Z84kMQsoqMIoQTH5yV14g34rb9BWrH+yPimt0SDth/0DL
Mz9dXDl4OSj0/QLrcVLHKyN8kgjl+VSMeOgRDs76JiumEezjBlHjKndN3KiCWZnDxzzsPDg8t7Ez
L9RQGn8CqqYRhtx7PhaQ/jL5kzl69fBk0wU09ofize/qtLAjqKvuiuJXlMi69cronZxc6M+RpSg+
D7Q8YgXAG7fNkP+F0aZ+rXXD1dLlx4oTio2n4Uyc8uatGUKcxZMGTJMKJS9QJYUN4u15zGoHH2E/
4nNcWKbhil6dQ+PyVCi5Ml/BVONDoWGrqMj1WKhq3molqrfKPsdTTN5LuH061Sp4iKTSyO3bJRpS
4uJ5d8tGDfdKJVX8Q4lCJUEKkOePOLZ3Hqf8u9jBeE0hlZ039oMkfEDOFBWlxLHsWuaDrCbXBi3U
1uZ/V22Z4p0bApHmgJ9rdZMv5s5LGoZzWgxbnRLwpJzDWA9x3vv7jo7wKPXwMVEL1MTu/7hiSYzE
PBQeg/pBzdY6OjVmZI5OU+/WX9CPnu/KH0aXm0ebjm+2Ko43i4Y31A7VKaiMdjA8Axmvly5Kds6h
BSsXA2NxIssUgl5VhvG3KQHoSpBlcbU8F+PyfY9r2UNIOgcK+IH4CaeQr20EjUXKzB6aL31Q6phl
32LiNUVd/cRqVLyB4qmhZZ1CTUlyss8OP2q7uxg0kFi/xtpMNUibV3/1061bzNHbWtGmulZrti8c
OGsKCBrEJSJZYrql1/3jo85NhaVsNNmQPWb4T+mHpxrTsQPx/oEg70iHSY4TGbosvwoxmAFUfMHn
UnxuIK9LXaBcywqe2JirsinmS3e+P8oVgibwIuDEZH6sGOgXI7kNLtHjyGvgCl7mehasVP/e3uIy
bKIT0qdaJj+NtVZgY6aHsZvGrikK9JhMFBpHEw6kXhRbPlLVB1wZ/Jg9IbCS6Sz25SuL9on/CxNB
edfzV3x0HZqacj3VavntDJ9o0qCohXN3tDVl7NqGCVSCe+Iu/USWK1KMtaji8YJhLxi1+RIwms/b
Uv8Sngezf/DrsMdkma37YrN2DKcpyDGy3cdLaK5FC4VRiEcSKIY8ohLQN3UgNUiDbTrQcMoRkgH6
6Gr7/DMyDijyHDXAMH3ZEFAAfLTdoMKAAV350mJD2TyQ8UKUv9k8RiIA7u+RWfn0DtNSkeDglklR
geQCBf8Jz/P3UCkIAC1TOKzVXitj64ApM3vChOOaoDzeZIAOi45fCYHOz/PoJ632QA/5vTZ5CpHn
YXu3ZZuSH98QTdkW1P2oBmfEvIXU7ZZ04hcU3vV6JV8yixBdTxCoE+4S7BysUF6FJTCOpZi8VzcU
eEYbMyfUMRQh9UVDuKxlYcsb+JISp0lR38XRn27KtMtfGs0lgIZNms/7JD/yG4xskskk+Hs3ALrC
mjUCKcaZsT3zRTwOjqZlMLvY+QSKwhL3mYi8h9b+X9tauI/JxUmYMAllfybDuEGdBrVvvsJ+zR+n
/oPZWcBUYhYIfRfY/S/x+2nCtuArhplqvZLN+uHlX7p7NheKQMYrKD5Gq3osVtHu2CI9ou4RzLsr
WCMG5etFG5qDq02PbgOFK4SKXOWRvZ9UtA+ePhoTAOSS5QvMqylI0fHAcdsepfVMbJ3tHrDqnuMq
GcQZ+R7gqz8dVd2wN+Q5UR/2yC/6mSQzO3KqNo+2YlT9qLxu+J/fKP/CAPDU7WnHh38Y8NT8lBZl
Y5m2lDwmYlgun9rKCUFBcGdkD8i2OZAG4Vxrs5rbgKhZdWOz98gVABSbDFZEY6bXXFWCY+iQbOBi
iYEtuze2KlOiFi12o9KYWnuI9ZqrBGwinSKYNPbnnlRinzC3DjiYR59RWfXdATglcnJSZfyzCGaj
fYYep5S5z77y+iGrwqdB9MDri4fPjdMjIdHpEpkl5+a1GQ/drcidgTbou2WxL44R5ItVp8OQMlwB
xrLB1M49+WQwYhFs7i/NgIdjNvoogJbKWoUlRkpj0XLTVCcY9IQyh3f/Z0xLWpyqUpZRn6Kj7SQj
fTXZOHFYRxIh9UsxrtWlpEqlqvddMs0WX9AcjCHnIOqfPjc9k2P8XeZIU4RGD4W5BX4lwhtd1bhC
QTZOf7YPEOKOS7oMW9UD12mmo6houV5fDzgycZOT83gasRNXSju4dy3m0+rqnGQfFeZwV15sg6LV
GYJmKnI1bWpjK2ZOBLo8alUWA/Pwsa8DdMqKlD531wgid8Othj+yXkqa8FjP+Wo6Vpd9BQQu7/dx
jgAM46mzFLQCtgliKDuKdXrem6CgIWYc96LT+KNnX/tGKPdtVevUH9TQqq0yaSxomE/lIkeby9N8
WYpvZfUGzFqQm6Q2E2KG7B/8aLxZNVhhgu3D2qjc4mcWWvqr/vRBh0TbKT9HZQePzuuEomoz7soB
bhgB0q0+6tomUvCOjjFPBtexIm/3XQGiRTZ+IjO7PK5UrDhORtl7U0I7bQlFyX2hGJO9iERnBfie
hk41F5Svp7eoBpFuoWV8KcFDi4gmObmrW1Y6FITFch9LnhHoZhOcEuBXvwF2uFYvhWGfAt0N+OMd
1JG5rjQRVAQIY71fsOX6aoGfaHH1hFVQi1tgHipUaipl2RJibR000j7tnmhl86BZyW4rFZNalsUb
vdvTluseV7ztSNv3+dCan0quGA4gtPdgB0j3a2OmCifvW9ySGefMVB+T4Bl8ypyu8O5Z9Y0xWb2w
sTEYDMqHYV5ggIFgH3t9QUJwg3m/PDz3ePCl+JE7tAsDG1jeKuiVdqL6/XiXmnlM4A+35nqx9wV+
xtqnqkDO2WINv/7id0Uw2dvOoOyRAGrE59i84oPZXWWHCHi+Od+xirmmXlHXv9kA+rb9GPox4kUG
CF/rR9u6NExkCvZxN2QVsSjk00nZr7T6KtHU0ZpMa89AEXmnHLrZM4EXDmQm9lbCImBo+oqDCgR5
qMJC0zVPoz/xs82ZYnfdAVcw3QWWYhVrDWj/2dRbOxFfyXkwrHD0iFUIaemkguJ+IisGVtz1E3kQ
8UPmXHNVHO0ipijI27upKqUGQ3xGxmJYIqp12yWKh1fMsCAkd4ujC9OZEk+Ok8ufL1Fsel50qXoW
OeHHE9gP2LRhghZe8d63SmY2qvJHspc3HDBgunirse4iFxpR6i/c2NXe6/p4bsqLMJgxl1pXr40F
VuKbIp7fvcSNNI74eHZNfvmcPK8TZTFWGO7VHJHasaKe2MJD6F+Dax7HFjZMgHI8JXiJlHJaw5V7
AxgBjDLwRJDy6hYSRb/GzPZtDhmG76tQk37rhNchWGMp5ah8r0BhcpL90uaWdHbNRzZoQJOXPQh4
aQsQ75BpeVx/gQyHHDDb0fPUC2JxKTsd44nKZGZZGrs6qqjHLXEsrDq0qIPCgw5O3rxRCEszyOXB
J6jpFNgqCNOK9twZ8TSzDZMh0LQnUMjHkSl82vrSAqXGsAXA+5D6EkilLOxxpyUM3NVkWoyCCWD2
bimuyKpF/nev2ZJEBsA4s4FWx1YFFJPOW6cpnNwOMitL7f3O1anJl5J0THac/FDq2fYOpTOaruZm
jALVFeo+Fcdb/SSVprRC/mHWRv+6YjAkdOAO3hroTd8pTVHTVJvjFsjF6qYJmwxwwSF+XD1D/e0v
fbdZRoRWio9L4R0q6k9/L4QksPItiLP45tq9ZjlpoUfxSUkiR420dwVm19ZPVTDKXS+b6hRJwgDL
T1v6L4tz4oupwpsltg1g9GGl7MlRVReWKXMKTyFlia+UqECROL6rDiAj92oneTSoKoSfiuxbD8M1
n4cbefZQVkA6bn3ClCvpyDwft+MnDHHhZuE3otbwAI5rD58/9yK+noV+g899d5jk+bMhaZnx14CL
JfwoYpjFZ0FHr6OaovrPtco3/TV7end7xiX0UkWKgU7RfY4lbEPYVkf7A2sLrnD5QREGp/ZtJWte
SjGXLSNoMDALg9URKpAaPycgUoP1kPDLJMN7fbhPrP7SQCM6plmz+JjP69tKxMvB6KDG+KU/x8in
HUvQVLIk09YpQernBPIAmhaClm0kiLeJetHlNjF1+R1cekHhvek1yYpYoWOievmqVlRkAxBFISeY
rh+3SweR5SQOJT0DhrE4hutsj1XkOMav83KqBYreHDzD0OEfgjq4ptQqCGWDNJgDVrbQ6DwMORsx
yrnoPzFhIrZwdzN2jFbaqq8CBNTvIUxxrJ8CLJcadnfJje1EAOlPE4FHv5qAE9vh6TaH+2SbKYmw
EQST4C1qjQB7wruMY/QEoO3zHewnfGjJG7BvrpRiGQE9WYl23ELHVpmNj63HhEwmdaFsMfFE7/6r
fpd60r+YZ4WBKQ3hWmkjPGDKf373vlI3LCoeYreuQqI1XiBlXjknz71JssxaW6pHxs51rooS5EwF
1LV9laC/AaKLvpzl3XLMXkVosTwhqVcf+Fxwrw1RatDC0UjMuPP+LxdJ0qrSJxlPhsZrj5GVBJwD
QJFZOsFBArA5TnadDA9DIbesRZo6Sftc74b45h0Iodx5nuj+yMV4YIOKd524RqkYsHypwr1p3/lq
QOOZyp70jS8Q4J4hmSa5e+n85dgxpvDJKSFV9pIiNCXQwIXlc1WGTXKOkqCvaLsRl5gHGpHczfzJ
29U3fcLKbbuQbtuAf5I1SpJifQ5Ou37/SRJ1PL7hbJXClM8pLQGDXAjftE8jH5Ae3iNWfdkIyxqn
Ygu8hIUkqU6It/EV30+tufBI3m07EoWg0KT75CMeSg0+Qo/6E/hKKrGh3Etfm34bgBslX6XI1ADa
2OPTeNjaEAA9i+mgoMtDbDado9nccEkCeeenlui/MOAF1yKeK84uxG5FyDCMKHeidBcKr6y4AfY9
GujKSzvu6JlhGE1+8//upMMFg6ah9h+SIlvLHmO0FPaRR86Ugo7lynfrjmTCDU+jcgX7oy7oQQ0P
DGx9fNkeN+5UXUYondpw3/pdVMx11YbohmdNJ3YYh9BUcIFGDPcBzIK9i2JOPDchAdn7QrUdjozA
kjhsnawjS9yPqN6B53PpPiNfAzSEZG+U5bGiBXFx/4NYgAQqVyiP3ORX17NY8VZxaxlRl4a6M6lL
R+WiLCKAlJUuGQhoBxs4b2c8PWpoB5D+KR+HcbGbCIhjTWElw3dnKK7D5y8u9MFV9Q67ntODSCCL
BYRr7VIaRvKTaPC7eRIuu6rXShSFluH/tFX2ml8X/Z/H5SM/D6U8CsS2hvASftNO8CDoE333KLOH
rTOi4SDFm6Cl4DMQ6kmn79IclVApjja6xGZ7/LN8/1C0AHzRpPcYLA4l5gs9HGGaxeCF+i7Mcz4L
9u/b6it0uzmY/JMu9QMrzoNQdeEpLGiFkNgl7xqhOV2xLmT9uZtnaX2orpe8KPGvw5/XC15og8eA
DBO4PwLabjU4xkW+InVeKb/eakKSPI4SyWG9sJlH8EDQdIor28kxKV4xLwxega/Y0PgKhYTOWA5m
hF63RCgzh17D6tOft4ZZJGHuiKbUStFU6OcvpQ2mNnMgokRIksPFz44fDAcm9188KZPX4R7F/+85
LYIHExGh1f4JGfOga945Wde7i7lcyvUM+wmMlmCqUahVai48XiPy7HArzvXAPtuqAWMetDRSy3ao
RXbilPQBd7FRm1YW44L4dakPqLPSWhBWSCFM4SKL6cBeaIsbtZjYa0v/GgMZsWSKezMVAX3jtsbF
x1sDzSw9fQoP2jWzK6EGj1d/JIv/FZ0WPJ9lhYBaCsnGabI6XgNxF06NLC8uUwLSYeZRjW2+N8FW
0ZFoEsCxNWYbyx33MfrD/QHkOT0bNZqBMWQiCl+Soub/E2jbvvftUByxCS0uo6BxnPfXrUbf4q/Q
9qLgmwJp0oVdpJOD1lalX+HsYxdDnfFdT5xTFK1R66bSqwedDwbBJQbxDUfsQYt8Wbbw32kdILRi
BhPoaSgBaXkFwPHIzkpA+SxqjS/PXkWBZLFg16chZGClPJifLDotdmrOCv2Irjd7QVHewviIKfgw
V6z2hR9NXMmdCiOBfcs+zSJs45P40pt3RFmzMJwWV8OIz6PNcMe/8T4It+lno5O592OVQKhBcdQN
hIr6MFDaziT3egsiOByWYVcr/6CkKIe2xu48EXVEfUjKsYgAUvyXGGsNn/YXZdUx1pD9lMPEbXMp
aymJXj9o1EcXPyl9slMspdhftVndHJG2bTa5jPSOfgtkLHjzSPduckiYAyR7UXzAznI0lB3Wl8KE
Xk50svn9jm5KDE+TFzJ4tRBf7qhwz3vIYzpjGiujg34b0883oi8vsLX7WO7w9FR0UTQayImitnyA
pstq55wo0p1Jwqzfjg5uZjFzHai34mIeCdQWhA4rT4daoHAx6zUXi6mRz+2k4k3Qj43aDvs6Siv+
0sLdfxsWJqVArkYLHuFzixTaIKZEig4kheyzQhIkwEt+ape6oVznyzMg5trrb94IxJwxIf9ncWvJ
yZ5+nDrJDp60BdB6fL1BcE/CKp8hdeDg3E594UlqrDwarzL1PpETi/L7nofH/md6CG82jAXF7oP8
KdimeLDf9QHqMpvWSRoi1w4CF0+KYPEtNvy/jYWiuU/3o8KupUgbzGWTCyP5vswfhewDF65uQZDI
kNdstJunuaWT6qNXdVHcNyezLyLJ/+yU/wMRYlvDveEyf4HDokybzTEOhBQyTUlcKpowBbBKnzru
f9mAKXYrAJUnPLLe/wvOxiL0nNkFhdYDfJwixP++HEO5tOt2F2hN9lnSCI8Ewxl3xwAxoQ+dAb4Q
zWmz6uQtasz1PmpZ9treS2f6QX4Hw9T6Cqu9D5x84Y0vYQXj/XF4matecSvmQ4/fgzWVPSR22bVP
kwOK1E8W7IcaKwW2FLfwYgJRT/G9ZXzNadKDAmL+pCTjzIzQQO73a9LYCGzfTfUlrU2Zw6I9uBR3
mOrPA31XckXnlSTkCO5tKL1w5D/6gcgRTUt2Nb6bVJaUS7qZIg2leKAzfuS7eWYJjQYL5smKTfQU
CQA4JPnMcNqefbpYOvGfAjKBxcjvZCtaZW+xkylrdw+zKEP1brHH2toCJ9OQPgU0LQdBIROu+zLD
UvApuJ8BQNcQH6nr/l7bjbMbcxps7udklXBzpNB3qlMG1SUrn/xcg2Z0ElE1C4zkWEwi0qOSgmGc
9I8TtMIrEl8zRQtZgZVniNs5daU8WmXrr3uGIVXBbF19ZaCOX8mVJMoiovOvaiv7r628rWJli7PI
uoI2QorhipMW2m/zaxoPF0gmTbFLpE0S4VpKQWV1Gs1E8k3/F1a/GEYYwSmSP00B92otkSGa9JYN
uNB2vl8XwvMHv8DPHHqXCcWvJWORMF1JZc5G6Ug/ZfIUrhlPe861OiC4z/DtWABJ05JW5uTgW/ID
GmqFQm0J+aSaS5us0M68RziwFz/0LmKRw2AHLQLD27mp8WFAROWULEb/t1cfT5aH0aVkFqgWlzEs
sJ8WZI4ravNVnWu3u58/1v/jbB+0RDcN2rdkFpKR56KHa0Ah/ioAdf1UNwTFeyR15mYmBOpA0dHj
O3XWXmN7Yss7sE3YvInod5keqeo5IPeUjMMOIFBLvclbYGqs9GaiQXeWAGWS4zMxjakDNMpNya6V
wzLExFJSj753zm4R9Xyo/R1JZHBcoWLfu0tq652gGmYB0vo0H2mepR2dlEYCfByfplfswHGp8wLH
Or14McM6V/C7Ifb4UmdbwIXS00As0/W0nIXjcNUZoYlgK1NOXGxAs3tlzHnPIDw8HSAHaLbWrZJ5
AjQrjmDVzRwzeZJgB0B90Dz4/EqDAMqO1OUTjriLJi2l+BzX//IMjq3wO7+fuoZPUaqMZY39P4Nv
Qm/ZKMWhYIZPkEuah36MXNwbUGF+0ucoyk8sDQMRmcQ1klnFY419Aykc2hShc4x9D/3364Q37G84
sXLSjz4Dyv6KSrf5hYocnI0ENux1C9ZCQbJv5BEd6bzbvTmESRrH2iZhcFT6Cf0m6Og31wMh8OFZ
AnQpNh73y9qUwSyowRI04gCK3fev+sGxSUaKuJkXBpZDrkCVwo+Njkf/fuiH6UEt4PGy1mo9Qkbn
xrDhp59JD+VGzPdd6Us0thyfY/KVLS49aD/IiH2Xd8/0oy55ULF33DiHnWQWQjBC1falnPH57xGQ
gSZjKFOXmGPs87Hu0T+QBjhoNbcj7Syu8k01QnZ8hSf/aBDrD2DUPbw7gDIFYjzzxSpImthvFAPK
ZT8ECEydecWZzxt4DMQgxuMc0S/eROHIibq5//KbwqDOhrH/8RNsCUa+zDqxR0gD1tzUQlOPAwfe
rCcHPocUfYRMXhgtwrCpfwxzNK0DxCwxnmuxkNmpUGlWLHWogxAF6AucYpfxV2xDaN0aEh0T2FYa
e7UewVy/pkysWIBBk3sFvgWUzSRQP3nEc5/xpe8gCojaudINQ7HNALXQDIkmSgeDM+ZLkbxmytJM
TgVWoePEbzR+uEZjDjr46N4SePcreuPiTEsbKHlBegFMioRZRHF7HGHUbXB8WQystnzHYqRncg5g
QCv/8C2+JeBtCKv+MukdmsOjtKeywECfWZnLE1f9Zaz20glRgw4bVz4Rnxz02ppL9onVizCKfaD3
m7f7z3/Sx0MjtFny2CmFUAwQZRvIveCohD/MMs9YVrzMXn8kBvaqIAZrZRZ9noW/A5mqsMw4zuOb
jkj6GlVcRn76uxrLPoDdWxoiSXEta403PK34GrlQAvRFA/6mqmMxlm9AUVmZhbUg2uJgEimeTd4g
3flK8dYWHHC0JDDRO9BNYLGwbCBLumupHZ7tPjvR667p1o/YBa7vk8Mi+odClTKn8j27fOVgzWAk
amGssUhklqaM///IGumd2bfL4wbFIPJYDB+OkNaQmwiEKXTZh9Cc4uI3tlSunJ/N0PAfBr2zoRyN
teHP3lbv7t2Ymf5xBeWfgnv/zgvUQcH7jj3ebGwnl+pzrcy7QCHqrRhFG14IaysJquN2E85ugdcd
iA+H9aVXDZ8jms3X5pYplZTqr5cQqspac+i0EkQn5m/E976RH91Xeyn0la708RrdpktOtp0+JQw+
TneYnKj9EXC3+bekLGGoY4+M6nildE8ujfJBjO8c0gt1bjorghRdvrjl8EcA9Acx0Lux1nwxBryI
zk9BPvqOE1SATbKHp3Skahs8jUju9wKo+VwFI+OQ4Jf9F1iGDUVO1bbJp1QdpW9d4WinNHc2bub6
5vnCP5FhOcuNgJW3c4/rDszVrEUhkEaBgGj8SdxH8Hrqt+1+jq1YQGFPuo+ft2b2I4hBc3PJq3Df
ZOtuyGiybMP3RvvINBrmJAnG/QxRevymNCM/qT+yM7lHrlwLaXaP7+VYzOcwUcTdQSQfo8fAQmSa
Yu7YstCtp5iNuOdQ7hAojTj/g+NK23xJ0f8v6b9h+RCGQHMj/3bb4yeUraxj4yHeqnINMV6T2L+S
z44Ki1EVWZo7TyB4x+k6ybw6x1ElcIv16ZmZoLwqe51uAQVVT7+GlzWFPQwxgqzXBdkvVbheQBgQ
dq5rfJAT7loFFSukQ60//tapz9TffvQFiwxKe+FcZlrc1/GaPuwbeUwtFByVUjSTAy5Olu36G5LC
ckNPszByyy9bNs7C3XCdJ3mfNNLvJqJWhbZTZWmHEFEF8c7qvRlm97LyalbavziERjQRlnNRhNgD
NZIusesvOs1/4uqeIM5AVPsKWaMnR3G7I5PLUo3ID3GpL3H+v2mZhvDmuG6y/w25AEW+fgFn658Y
85Ajgzf8cH1o3YlrZSVqS1PVl0jWQKKLJHCLoVrJPqFVxQ3MeDWCUeqiuO7nWi2Y/+AiU5UbvrOT
SgcOKTZlskEJAhw3JRM/aM/aWSSim0fgVL9lvNazrGgUiIq+CVfOKSsCLLc4QxWbDSRnqsU9Yj97
KB9TQm1ORECsKeBURhl0SbSPzcHXoUbb/o6zPfJ+LXWHd3hp7q5UAqtBR3tqMWvCeFQtcO2HpcSi
GD4gbWFrooMmTvN37wOGxwJSAL/0g4+CubbYNvFLmN7HFzLItn5CEhfZftfoLyZgB/lbPzNxG7ZZ
b83UTcHaeKE/f0yxO3RVo63WVZUI8Tfddeos2Oy95sx7csDhiMi5MxYIB9aCwAyuE5+CejT1w+Mo
AeW8adc1aDBARwpjFmUtsejdSZXVX7um23Kx/gujJvSf3Mx2+3B/8Pt74b4xPWApb5gqC2n4s7Xf
uFOOZJGTPC6XLU+kHEMH0KVmV5QslbQ4lKaIx4MzhYR0DxfO1qxn3n0F1UC0WGkZPgabjIDJpvB7
OYDAm2Tg78CVLBiav2oCknnO1c7twCUBnpFAIYriJLbaJ+R6N2NRf+yzAXofT7kwr1xnJVDb8CwG
dHZ9DmiT4yDrMzSGqpWcfCfOfvIP78SABfPLFpurLK9ptHe0Y4oRQucZgSvr9dHUgrclqZpSwlD1
rmQKTY0zcL7n9sSFnWBFzAGEnRciU8zPX6Nu28RJuqBfipBZ6xku1uHe3KewydO6A1IgrBJrv9Ll
3ACAxeo0s5ZWbT+b4gRnAyGSEG9vMaXifWo15+L/bVRWEP4w/xZgRnyLdmfuAj2VhR1iqZ4/O6oZ
fcu0Xm/0zRPX0kqLIB/YlN79e/mXUXf/EXVXaQ4CdpSiRNUOSGw0g15UIItEi3kSEqfNq1u7kXmX
mLv1sg84qWlYr6EQXaJ9nBf8ALgiU7EhSTR0YkPwv8t0Mtedk7eSr5g4F4Am/JCDvuF0GqH6sVNY
ED8lgut3XelvXMAHsuOkCVzWedwl603+xJwB+SHRSO+76DrEuo62uTmsm0PeBwWSEWh23HGeTIbz
a8MlczfVCjYFV6yw8pR4fGT1enkkxRw1/eLr0klOCubkaO2oDbnTYQwCRiOrKTNgK1/j7Na+ya46
/D5zbIUNRclOxNxNBz1hs92C1EYkoYCw+RAqiZCEh8BW/Vk3bqQF7lqETbjARqhTZT1X23CoMB09
/s1jONMKI4gui4gWiD0pGzDUXNur613D1oKGsqoIQQpAVrPY8iWoQ9ZN8EyOpRlFFe/833sExCAt
dVzIHPbhbj6pbIrlpMCTr8jYFf3WpZUWPJGVj6N2slPC2NRow7oWv9UA2wuUiNLX8neh1wfgrEnC
QuLjr/croH0EIjleIroNtaf/CNEGJG8wGWW0EjlWz5GVGfSdHiMzDNWqpdSkM7mLvXi25zlRuKrR
uNPBja9jF6KQIKOcjfFd0B/MmwmMUyIV81T80TK66+CjV8gr9Y6WdcB4/RL47QwlpRz/qSsVzvGE
njb+TLFZU3lG9YBR+QSxPsZyaQKnHhsRVhlVVSArLygDhyXguxoVDFHt5/STfnEFxCSJr0wvtO3v
WnXzTrN4tSKd5TY9IRJwZ+6texjXgSF6L7HUzlmWUTk6DJqSgqWZIy0hEHh2Xcvv64LBalqqVPuh
eSXl4eYrYOxplD25ZgOONtiTcIRCuV2Y1wwdmKbx3WclBARDO24vqlm4KnRLleQ+Ml07haHO+uDp
EoTTm2xE5ge8h/QuHD6rXFOML6WyQd1YoJHJLUbl6Xo0d+C2qM9tBLQsn22x182CMNefCv1Bhlgo
M9dGGqzG4VCd1f/csbpruJ8eyrIS1caR48u9Cx01A34EJKlL1bd3C3zec5WGDS2a5tSi96geVfyK
njW1OPgViUiSfZUbx+131k62fprPr4fBfFOX9bPUNIjypxUeinqObR/iW37za8S3ZDX2gLFv+bX+
63X9ggfZxxZWI5RXZXCSTAWTBdWTQiuFOexBJOUSBQkbKF17jnfzFhDKpBtO9wf1PxMfJ8dcqAQd
5gVMeTHZxwePD9RpsnLoVmRhYnqpAIRJzHi8z1Yrurwaizh3EwEM8HX2Q9rDmFEJ6i8qbVpBQS9P
WKcW4Lz7CuL+oZ/XuP8b85hvIH/GruwoXtUpLhg/7WbDOANj2LdE2GzWykiekueij5wz2Wzl6HKe
DwGKg+FUr7DZvUvCefcfleWGpM/kwfCjmpGklWnMLO3XC0hktj+b7bdS+80Jmrb9klHpdOGB/8vO
8EHhL7BmyuUIvQSUJy0vGJ/fMfsLiqqlmdvXZW3zhoKv5vb3vVY3Qsm+lQjRDQKSrRzac+lt2GB5
Vg6LWuVitL8VQ8oqGZbJvpcsmoYmMV98oWyGiUaLpHRH6vbwSTX82t/0evx+Fk/t0e+htitXn5rm
fAUmMjk17QGaotFw+fJsJRWW6iLrE7qZmCfxw0PXtjuoi27T3btTBxym7aBgVAm1bJCDhxb/xqtI
vmHvoRAkf2hKuh0ssu17TSUZI9iuY+GGd6Q+HYOrvpMv06/GXoNHLvk+/jC1mnHF1GNcLVvPDz62
RCGS5/ZwzxNL9ZLdbuZw5IGbbjtD57S8TPLajhEZjqy/Jvn7bBdEdVk8okFhqOq/BpsVjwDxH0Ml
1Kzq+N4dZoQnqc546n8X8jp7OVGaUDSuBr6MGnn3inOCzmETDg54bOlyYhCIp6eKssfhuP1NPiB8
kGbghnpFN9nLKBcrlzHDsX1/ZFmAePnvTU8n0qxJjguGJsXhjPeRBgwtDIePUnrri8QPRHUH6NzL
UmsWWeImyEaCn1Jgps+7kEhLfXURRQN3k/8UijnR92FcQpfJFPU1HfJ2i6cVDbPMPn2ngS83NsRS
ZAgpsk7VPfrC5cHjZKiIchM/bgUsx0EBNIyQD3PHrjKHvDXVew7LMrxoxn+lAyXNoyJR9/sDwi1Z
4DpjRyvPUJMD93SJ2N9plGQAr06KgaKp5N4X039ZqSUbbRrQyrFZN9u/UQXmY7ZVXd3m3frFU39+
mwsTiN0ImEFJyIXt2A9rtMk0FnjrYtdRl2C0QX1ozypycI7T1tZodVx/eWYFIjwDXdwviUbKNPAR
fpQT25q+rji2WaxaMo37Xo3f66eakw900qPTeugaCk5/3IUPSPFxUZ6wG1qLPdRCckd/0OVJ/jHv
1UrBR/rGllVom2PnWYN2k8nrCLaiv3tQjHnNs4gcCQE1ylXYRmNcHDsJGImSy6vUko4HhnMLxBzn
9L8eh7mTkUPeC+xO1uMBTEshSFEH+HttmK+WcnzjfOVDrjOnjAITGYSBj4DhUp/F81YKvFoehuHy
9dZdR1ErkDRDOLqy3eKj44exgkJUhIlk8EONKwGL0frtYfk1ZPsjSzoj2JGhWpglDbPvg+hbQCgf
5RmdJiONVc+7mdzCAv/nH6jgB8BDgZ/gmsrckIDcFqdDQtfb5AnLZuJGUlhFezh/JJLEOlq/1P0J
AXWgqVsvkz9A6wAYnF5Sn3z7ZOvO77e6eWr1wqjduVfv+V798/IhH30pvoEy0DymWgQt7yL8H1m3
oNHpF/vECqIE/c5Wgtr/1V28uMQXntE0qzEgeVJxZuky3Yknm8rWgjPGTiY+3C/7b+KfjxMQbRjQ
5Arp6pJluzBxGLxTrr6CMGfIQjdo9gp/nTPsjSoqN4g/BANQcAUteF/oooi8kcx7Q/33dx0QNOLM
9ZOpAr3zuYB8yyJBOXZqYKHT+it2ZdZg/FFmiDUk2eu7EjAET0Qb2vQJ5FmsD/TdAgwUVuLr7Hsx
jPjC0h6KopaasVWrlG7LhhskVLmXdaiIGks1GKiYBdJiBTfutxdg5pqltfC+dgCaSZF8ABU80l4e
XIfkGDAhYHbzNf4pMa/IF6MU750VWWacVmBC8BqCP/HJgt0tvtMaDtxAGQhm5bjiglCvHNhxgq7f
UscSco1nJgaA8X4pE7IQuS4czlffLk9N9pfo2iCttcsrY8gcc1NQnOilsclnFvG+HiGnvXQ1FVIS
wQB28InqOp7dOK2JFR9wS3NHnP2dU3dWgvRRyj8JnzFeiy34idyGYxrd10IAniIfx0zPk6BlpbCD
b7f9wGy93eNL+lv9FeSxCMPEl9sKLYvg8Vcxy4lieAREDhibvgbQQ9A286dwG/F74CxqmFGMAavm
+NEjSLML4Qkh2Dnq04XnQIqTVq5XGghvn5kEMz1KLmqu/H0RxmfCmhjCUwHU0PyI9bLDD/nQIM24
zY/JNTX4FcL2HhK+fsT4KLUEIrHvJLqU/JDMnYNkcfGZyQjGmeAlwt2FMakfJZGhr5iyzBwmNF0i
paJ1CsIXu0atjVMyNBgoBg+uohytwA65WvV35ui8c2npCYL6tI2EVCohhl2QuYaThp6a8Ai+zHpK
wkk3VqhRVsrWnOAisySn3eNy+TbiA+MHeNVStzPfzr9z2g2yAPUhwftN67Rl2EXw+TJPvc4COTYX
Dl6g9ubHp613seUSFMDyGHhq2hkn051B4i4rvyz8vPD/D2JiCgaaAj8rHG7dbnwZLBKLSZQpm1n7
BReIw8O1s9I+pg2L0FzApGW76XtTG9Cy/TN9wxGGUibutoTnyY3k07dqSDKwZFw610ZsbcW1OX90
7f5HbI0Xbfoc8JJZkNM7BA5K42V3Xw6LcB2acAEfu/xMt36zDB8Q/AHL1lFk/34fnkogeTgREiC1
VhuqPJ8iigFK46tU3inEfYu9kgqXs/vinjvidLCrkouFazmRjT0jDLYSrUZpWats4rn4PK754TuG
hzkyMmasOWG9MjtGFrQPUfGqrRRqLwBvhRBJuInWYgsvGZ3NPKqejtugDmGB31NMuxTmMEQebzuH
yYxifTApVvRXdGrEzTKKZvXanskbOjv9W4JNDxaJsP3pLFFa9lkJ39/BEa3Q4X4O5Nt/nomdlZXU
ACpMoGGGy3tc+z1Rrur2woxQua7eyDbehFCQmscR8+ApvXHGTagPr4C7/NuE0NPKTbk7ShjhF6gX
l/U4NiHZ25CRae80NEGHEkINO46Cw6WXIU4Nv8hqVxRYEkRiMlgr52CG5MddIeK0LhY/2/Odagu5
W12Ldozi9d5XSEzobHGH9Bb2XJjAr4OF/MrJd1YL4lo0Dq6Z9q/gw4La0huFEOvUhnh/CTSi3a78
D3wZCY586aBDe39QPHw/vdOSw01dOgs65R1121HnGBizewZ0juiGle/gRIHhVRPoL6rVTwtgm1PB
RSb1nFCFBDeWkdFkgIENSsH1/M3/IFleBzan6n+jEuqoKmYIZy/QvaVyeIBeheZKg7Empt7erY/y
mHNY8J+h6FB4mzePWgjYuanYeYe+ZIkEKMrtGu+frJJ7XIQ82rdcJzNDU2VhRQKCcYMjqckXA3PM
nyzLZscEm3D3T19oLrOibbAUYOyxrfpUDrkVRNanbxsnIe5Ybx0ebTOXbTYoVQaBD+G4tNrL76SE
EH9UkLVIhxTSdiMqsgbjx7LL833cZHJzrhZxDjb6jsKpYAIKjz8r1M99sLn7hjaArCPVS34kEGrP
O+dVonR+kOdX/LkhxJd4GvSmUJr859otkP0m23tny4y4YAWmhdda6g9Rh4W5nKLM0qIoQnL1gdGN
xPVpPteCUaQkPrJH5q0/nJ2z/1Spa8tK8VlRgJ31RRbYbEl24/ATyzDka8ODq6RMYUpLrEvr/Z25
92wP1gRLF+2Gf7tmOhszodq0wVt5H3n/5B4cjTBSfqMk3oII0grhaKfokPGWk/V1Flu1ueNK8WA+
WTBb4uAE/m7w9MJ5S7kSTDCX5287Qf3wbU3aylU/5NNa3ZM406Qz8VZRrBB574XZkSqMI9Tt4bcs
UHPyYOPLxULPMxQrHsy5IgGzXIHDjXEXigbKiUPLqP4RTALJtvEW++FR/sP2zRkNLIjGG4Fe0No9
Jj5NiAWk1LzjIxWnt4jpXKqLZQyomoiHAeN3E6qMlJMVfp3f1XzXvv9CffCcSU1wG9AqSfje8E84
kH6NN48RKztyuMMfzQ1wcOUFKxOomMEOKllUOHYd+y5D36qyVGS8jwdUJK+CDFdJ+ARIaPmTHViC
Z8DhBe1leZt4tx7GY3pmeoHcLrbjeffa7Rw9dJZArR7vq7D+R9IR9J67Rc417BpmxCyL1eYhC0en
zgVAQWdG0fSndL8/r897G6B02FyWOOcVRQ50bClmMvLC7HeqNMOrxVnZRl/0y6/6Sv0jB50emFLJ
uQold8AvJHSzhLbwsKmUjNp3+KuMMbA2T5OV1bfCxaQpdW9puUMmfnHWYytBwTFEMbG4ghbYaDaf
3v1Y+X9mJeLud3V1RHHxVzpiUxd1DF8JTUiCubmftFSLhuQ1cEdkplhaJLSRRWHN0dA4+HH3n5kW
sXA1WdYtcW2Gwpg9tFNP0x9xK4fTALcBmDkTCak5nongu8TBQ1C2tPS7ResxaLaDU4ncvM6cIwtA
EiUZbFbS0/S3Sj4xJoZiic5bg+dXaTnnFy8AO1NJzh6v24FE8304Q7BHZgMZHvfc/BDNx6Z2ukqf
MY8v0WskLFT7C7aOeMDgeOhoHNAlK3V3bbRDTreSndw5cKEJ4QoKF417oxghl4t9Hwpb5Fnde6Dc
Q/ei83ePReGXMDO5LtE6HQzFQ5n0zjy1uLZupQp0Z+JZEAixV1lV7ZaPyQgROSmZgyX8te63lDly
vfKcpxtPigvcIl3dlNNZno3rnNui4vmOvKHmjWYI/CpLzGRDmXij0enaWI1hmWhz+QkhRpZEbXAR
MXFEmo6UivjG4PNAjjoZED+I6fIgXLk2crNwKFpr5qA4BboBAZm6stJ3Ej8yKrn0a6156ezUB9+w
dXY1r/LXuWSSXEsT+7e3CwkqkmSq9RbtgxjwpRrgMU5M9ATcAJQQaG0rNKZf9PJ+L4v32+eOT9Ac
RLqg3RypkKV+w+JfUxVesJJZQzlj5fAQ8o89wS8I+u2C1AXOwe00tQ6OS8TXr2Wy3E/Rvyufek7t
4vPdly3ROT7xj6ye2RbLVK3M8VO+FE1q4eW/WFMJS15qomuKsG9VN9reAswIsQaKGRAWbIhzbGPt
9yKG4/EJia8zL15G5QXXsw1e5F4YCT8Hypp+NI+Vvfa2O8u52/kRoOBqtNvsx8ZmE24IlMybL920
/lFxZsT7LM1wb2C0M33x/nntg+U/rRZ5laepsi+h9BiziPK4a4npLOVh0DUmpIgsu/2xRmZJPLt9
cCN8V6ysh8bb4pTJn6qGYvJd83HqahmdIqTE/EwN3//vo7TtPgWzW3zQ9aCDnejvdsEAsrDs5Lmw
Nywq4Qu9777KztCB7klt/nnnSPBVEoUUybMWfbumZM8+MXZuHE2x6+Yii6htZoAsAMdpgSB7zQjO
cQSB+rBs0nxbGfIC4ki3rEDDxN3GZGwLFeWRJsHnIj0PaHrDLmy6T5EojjVygCaF/ZnWRjWfi28T
9Ml1G8WZLJKc/92rRJNncEfbCdcWvJS4jgkSq5K+XducKMRKGv6pMJvQSUKe4loWrBz+UMDXYsH+
zYW0W5oSsbNvbz3of9Ez2a3cFsT5NAiBSzsUX0g1vjpImjgo4Y/AGfYs2xUk7Tu6qhO4gwFl2K06
o7vtd4cpiQJSpYu3l04cRkLsiAPwx5WSGlmRdehgojEtxS/MCtXzcYTv1USAxtb0xZdAOLi+I3Tf
F6sJSRLxcBaD9+1XhVhKHd6oEUKYYLtubHu24C9t/DC/dPUPnKVfeNxvAeb9n/G0UKGMp6CO6uiQ
2mWzPfDbkXA8OccHzkUOAPricm8Sn78Yd+7cVHvDi4wUW/ZRoEZwyauUQoU7W7q3zdkoz67vQH/i
UQAZkuSHj5JoOieCai/vDVTc3ytFG3lLyNK9hjBlNbHyF2vgMTamOcJbvNOVVDOCKilia/yc22hh
YzgAnMn2/6DGGH/BZ47G05gfKiNqmxadhxYKmrUEHch7bjreyGBdP+AJKLlfvfEIpcm+r2BEXjoz
f2cxGl2gqjluhcfaRtIWcDo0TGEsjc+46PVPtIJQ3wINRr4NIIKkGctxExgvikWXcJle+9wOMmJY
6XvrfVKYyVj1f9Bo+tvAQBGlTOV6lXZiHE9g5RlukT1BnsMe/ltqrAfNten6Z42BKw8swdxf9BEf
RWkC/P8SCp4vQOSpWkb0nOsQejpKlUNte/s2WO1Frmtr89tJPYCwsqb+iWD7AerkjRnfn0S5ahJS
rNK7b1DJVmw+jvveq99LSHss+VXpoH9Yk+IA8WXS8yk3STL69vWGQDkD6/cYyqfiZr57BsxWBJVQ
rHsC/kWeOB+gXdxJ8lGqDtRjmLbX//XY6FprubDfIGLMTBGm+h+Jrj5mZp9lNIPM54ShtESD+ZfI
YwDVIAQg0ZE5MTR2SPavuUfN7nMpiELHy6EKih5LQ8vfBmN49WqzI7cS07erTKUQvasHHyrbWSr3
r/xD5VU2lz/ZVtPuQI31vNmxAwuO0xkGe/K0v0vOD97YxxInBL9UVwWUACScxD6qCJZ5gWDz408I
vgQ4/Dla9Oh6obWkKdzSeTqbhNFGld+26bU5rFWoTnqLWXO0pMZNC11ekF/CkP4SgKsTizmAwLZg
dDnHAbwZzkI1Xq0fNMXDAdhtou57RDj9GGkf1ZlpOa6EBXb5VziL29ueq8ZuyLYHt0b1a/AslCVh
Wbe7NwU76FPIkaN7OINfLki4kHZ/XLWjkv5vvly5kVdjqzsLwd4/78jaNfatZClpAycbCPzT8CYW
td6xHodbEQObIyumaI2KqhzLF8EsSq+wamZlssriVaVFS8Z3Z8cENX70Ib/hQDj3700J21LjL1UN
XNhFUqeK24omQTjO9CrxleQFf8S3zln2k/HJtn/X9ccJwv5xWtO+fRCgCTsU4quw5EBsAS+YM5V/
/Jm2WbLmb6X09Kls5/g6ldRE01KNXA9IHM5AUOCp3QNFtz1mePNfPbZe2uc3GgqfsBol19oAFtsq
E9uuxuMhaQTR2rIDLMWkA2hL15YQ1OwOP2sZqVCCg6ikV7jTF8IjJ2CFgZX7r4DyrlXBzNK7b+Lr
nhFuLD1a/9hZuKkLA6eHpkKcPnurLFkvRZYed+WzTs+N8tQ9noonuiMZp8IVLJK1Pv7zxjLuZRkk
TlY21QZM9FlIvm1ggFuR8XI275bFiH+GdWQtQCBVNKKHvx2B+MSc6MX00lnnXa9TOnAt49Vdhw6V
7CimbDRk/BE/tXxleswHDydySmT2RkQzco64PKfB+B42i75XglRMixpNAIhBzdRpWNbw/laaTqAv
0hIzPNauNV/XJNqCz8CNMsx/Fgh5RT+Uq7kfOR93H8Tq1oVakjOPQPXKOrQnKKsSzj37YRrxxJdQ
ofxedKEUticp9LGoxOWLYXPg/1jByn3+hgZzzLGg6XfXoVk8Bl6d6rBy47IixHLiqrlxDe9OzIBX
C8VkXSBGpkyh6NWlwja6m3LKrK7yyukvlAyfPFX4P8pwVSZTvmiBuGy2b0KScOb50LQtain9uUMS
5yA3D7C1MIq5hUL5JrZO+tn4p9s6vSrD4OeLoo65sRpcuQ3t7cpMTLS8ISOgAOAL00LfYYj+F78k
Y/NhcLBhNjLQzHz44fGt965BLUBWwSX/8dEEpxQnruCkoG1bD4JnV37NFjwILR6ecyQC8GeGPquC
P5HIe0i7zo1xRm6QPAxVxeLpltneNDidz2SXifHzeon2InhvJqJNDdVXQYN9WflZZZVRbwKPNbL7
oUdP1giBeu1jE6ME54JGQcBI5W4MzaOYI/bs5MB3PfWfetIn40OxVwjfBTW5VZ/HcIoX1cyuyaFD
+ZZ5cCio+JoyTRYsADfBOkRGIjwDO1gHeetAW1ZFITp8XSqqN/4d9Ofla9TgsI476e9lH8LfPqOz
LTBQAE+EenkUEdCWfsys8oLjJY6KfGwFbcFGaSVBrTlIfQEHbHv47BgrR3qzVQZs4WqXnjsdaIpz
6ZecnyEZF5v0GGZuPlHGIH+/PD85lifkw2bfXF/dur5hc4rKceAAfv3jQ64AaO9R0j9K2TC3ynaY
yU85apt5wYD+SA0hPEQPId2RZK5/Io+0FEAO/75Lq+vtdshuAgZFnEQKK8NJa7jS0Zx8TlH/7F4K
VTuMf9GKxjisdTDr4DsBa6J5t/rNgKChDb/RO7wNpX2FUQCMaw+U55tD6V6oE6wZUnhCrTZfTvVA
W337pbbWIYptobmj/L+CLvfqj+CJ25/HmqrSCqMH0nelsa0IB0+km4RcK0COBkYBlF7VCdVfQsrN
jmt1XiQVADP5h3K7OTj6UZ/tV/BAjUyYkI0qnLMVGXr1n4m9Mith5SiSJc6CxHPxr775X7b65Fur
pE+lYUHj72+naxAVYHJOjvd+CORJCiM+JVbniV9ftHJBCBRTPq2dbY0Hmtz8k5GFHWZzjVapDHmF
5yuwMrsZ3yY7S97/CzeroN6NMOhO6BZoSt6OMF3HySuGyYUIPsoRtNd2h9qx/OXT/yY5e6Nm9OI+
DNTAF1CVFckwAHchPfGyYjv7XYtvy2eAROIOu5q7fnwQ/CYYUcq8lwc7rHGKRIfvRh0a6E+BAD03
1x9ZNSStY1PS3XaNQPbPB/f8DiMctblaKT/0r0w29o6Rdyh+/O4hexCAgZpfxQkaDBEVeSvdxJ1U
s8EEH6wpzXbSVrbSB4/knG+xu7oSn/9R2dBf6Z8j/Ewyh5flRm0DkZ+0/7gyGFfue8E6+ngwVCXu
G01iG+ujNCfm04OpjAkNJy1jVTj40qer2u286bpNSiVmoyRxbFLHYX5jdlQqMozg80wtQzF9yy0M
BPIxeAGRhEZzBFDpI8HsEyYQ+kyXyjHRKSlZaS6+YTNJhPo7UguyETIDHNSBfytkMdFWwjuV3190
qBDfR9ooMICEPyD6U5or5KmxlIjOB2orJJvykm3LzziDlqbcZdxphHvR/gj3httfo7t4LC2lVSYR
jVCmoQvf0fTW/wPiWvwksJBy0K5yxETpw0WrlQcq/aI0NESrWExo1Dv5YA+D7T01NRTr8mJeyI40
8DfCX0SAm/vqF1rx7zmTdUrWfNWG9wgAIlRx1wcUDfvxQaF0RHmam+tmeEh9E1B+VjY1VxjVIyA5
2WRw4XS5gSniNvEVTV36yosPxJEabSOHeShlCLwVmrZ7Yy7/LTRoFnWKjN+hRUmSk7ejMy6HdQOh
Ta3HTc8ejc/K8O3OgPPqhJ/hCoNJa6/quJ2xCrFJkPHub2My33xbgvTNi3KqKav2NqONdEi/tcu/
hK+0VzhM30rsGPIV6f3mH5BsDz+a5bwhJiURXc4QBQK/hHX5+e2GI8AIgn1AVoAr9WCog8qNuc2p
HXbUbvfF/B6T5QDG10YHACmde1jIGQPyCqozUMm5702wj5X3ZkdJlLdgxJ96D31twXMvFUYi/h35
5CcFVx9rgGNCcsmfpXBvR+Njl30Jw/lOeU8KiBFL36LINupbtiGCZaNDpdfzt29fARf5d2iCoScv
O5gXEL1xndwoFwKE+yJ//xz7/n/jfXTlviWoMPBx/9wevy55uyOeSQBEtvFE0wjnMc7qP8nPY8Bz
uiUuK9h4skMVG9g4iR/A7RiA1wYKVxAsPjvkMzNTZJBR5pXzwC7K4mOE58wOJVzZbi/aWwFRlijM
SJvG+TIoiUYjoTI4y31mhz642vyXL18cg+VyHgbonh0eTO2MsHpGcwdvnx4RGFJFlVEOzgiPRIsx
Jg6KqfbW7aEsEwyG+w7WqgklawHlYLUoyrFGEwJ4nu/j9f9IOkKMLel+N8knIjNHg0DydgvNTjS7
/CyamDWbJI8z9K5Iy7K8NlYg7aLBnlGx69LOwYjGnwXcMmcgyjGDJEq83FecObmyk4OpCg08ef8x
XwNT+B63PB9A4BiyP9LCAYby6+C0x4ljkOIL6fchJzOCZajWncAUL2ffJllKZtopkDV6/GWvARax
RUyCQE2URdUBczNh2VrQf9Tr1hq4mcXkxLUSBCtcY+jTFDdPSmstMKoz/fNUlDWgruzJIKYCuwWH
qR+Qi7HjQD/WGh0YSEl+ens9ekmEVr8xp63gK1J0bE5pcTAsPvE6KPSp9cle9u4aCUah2JdXFrMp
CAJ7YKvHN7cI2VdFBfTbPsRVCk4SCaYLs0XtbL42JFmbJ59mKN3Ddql230CmJK2Oewe72dwDFYUS
iQVhug1kSpJ28krpWFYxsz1l1q8Lk8pvHABSS8MzMrV75eGUiHTqlivD7F8mDFTtyHWoTWfpAHav
cieMHVooOtXkhCSbBAwFGz2keHcnmTIn5eHT7A0xqCGmB4QqxhlpSLr8LAU367kaR0UAW/kqaZV1
6WywLtvNRnKyQSwc7gPth8JMzvJYIuOm6VmGVxEGh8vk25ADnp8SgFEJSwYpWKZ7ikTFjKz2LtWd
JFyPGXYPQnJdJGZ0SntBjcU/scPuQguQDtqDbMNWteJ64g99qoZgDHUwG9kUDW/GsebV+E/zEo2l
Sy7VloA7eoIiKXoKQFNUvWg8fxjY7mgFX7TNQ6eDeJXhJWRbGh6+0TVVmObcxbRrFQ67rpSVf/0B
GF4PZUw+2k0CFr4T3UiauCFHxxXoKuB5OvhrLlbO1UuWvPpzfND42uB2U6EuULgJ/4h0lUZqnlsd
A7d+qzfPQ0lDdJLofspKT6mSeZmGkil7S3ctHxtWUnSfmbiqdzRwNubJILO41W/pu1C9yDS51UJa
q/w53c7aipLzHU13NFF6TK8EixHmwE+tAfD7rQdd7yQwAlP2GWgRDoj0K+h6Ukik6xcgmngFSQ04
dB9err+7fbFOMi6E0HL2svBt8Wayora2aqVub0Ckd/VYi7aJDos08ZRdQuFiTsyj/EMnve4WpY63
oiGR1EUxx0j9qEfyNmm1g2cWTBMkq0xLqz8fjZYcuvdCZ808Bbjr627kiYbVDXNK1ono4DjZI+V/
NqatuTtFMfDfR3di83wKw3l+NAZpluJlBEKGwq54i9MD7r04REFK6GBTYN4UBVZkQ54ejHBFJdaw
S0tk6vsUm8XhH/0qiEEu/tjv6LIeLMbYqY8W1k34tR39ZCRinrnIbYaiqfEnOmLs5eWxH9jnbN5K
SCteu6a4yXKwboX9WktCpXXUT+plqIAXKfEjMfz78gOaHl+dvIybfkUm7PUarN1/AxaKkPEVE50u
jZkstCUkyG3/AJ6zrRak86denTkTaN27O09B0WtsFK0tXlXkhZg32IKWeO6Ssl6d2YtOVZglKrUx
X5Vsqefigp1kx1hnRFL40bggHIE/6Ys1WvqMX68wHggcAL3OhdIeiNJj16VbMRPw1nINgHzLpiCr
NaSsKJbIwi97AXgvdI57jt1K/qIFPBdmWA4Z5o9QO+ocvbj3BEQpaZiWhQrAd8GYRwi6CXPbYYBb
2t3CkGnVEkH4UOSXid6bVeU3QstykI1TKkrUdgpNbLMurxACpNxHJiYcKrkhK+BUQ9V0AjK44LNe
asi5NqX+UxEa2O3nwWjDFRRqO4bzivafxtCbrQEgTTzWSsruL051scDJL7VPBIocvhUicbMVK8ie
oX//PddKwbbNeqJNvmG9oEWw+BWzVvzbwbq84PKD9OjdTbsu3zAtyr1hGXk3eBMyqZOI6PN9xg5X
ekmsTaAeZZ9MfgEq9wFTDGe7qe1kVMYiQXWe2La+7uftxG0P0mVxftd4mwl6wxCCtDl1uaNo41QV
MyCcycJIXMtyq22mJQsRhWwvhdGJpZEQGxYAN1ElkLXq881Yd6F/fFeU6M+plPFMp5y0xn07Nx9m
/D6JSDRoKBuqrfeh2stUYL1xcWIjjWxiThJHvEpcUJsK+jC7/NvhvcDNmh249mRusxwpQ7YBcplz
AG0Uw90tSDCAHQHBHWbrhTuu6x6lFTeULpxrOQsxq6CpX+EOeJ9DpW6aHRFSlwl1YTUbq9fNfFdt
9f86CTDonU+W1Il/Y8o7Jtqu1QSu8XCTPx9UZAmkQlHSjHjEjac/sgawO4K8KQbwaaRbps2RZN+s
cShylqXCY/+jAgPWQHSdW5f+5r/MHFj6OBnCrUKzGemc0EQEYSX/JqBZX8lmW/c3QQvJnGXpb+xi
edIj+H38RI2NuFRuh+Z/AIi6ogIcOuD3n0mgwu/5ryKT9yi+30+cqRNFgpOKvhBjVyBaUZcT51uS
xCn2QI/Ce5azGXH66zGOt1lVQ67+/JwcETtNikK+XeCwxi4iTIdab1VZZHkCuB6b014GrcDBLlgz
TXQD6l6TIONTsOqO4hGZRrs0QLkBlouJ8my2ShO1+u0tUX9xfAbnpQ3oxqGYvMtBqSy1A0EWVghZ
4Um1PPYSnpKom25I6px8lg1hyI1P0RnbZgP9uTV+q0BtV/BiCaCje732hzneoztBCKMcgVM2wxy+
tm78H9ESB62/XjT4KS001WzPb1N7PLktXSgqApnbqQ5GRUpSf+dp/6EWMffp1UEuOBB1u/uDn/ck
0ATAzkBQ/bjDaIQATTt/DiCTGU8S4b2DKyIzr3Be/klYQcnFI8aoXdK/xn1sfgbdDecQ0VflkZ1G
u427OLtXw61SwmD2lJBFZS7Op/BNKhMOvHPMEC9lg4J1QJJdstcC6Ypo0FzZpDpt1xo6/lpqhCZa
8Qk4mmO2c5FKUDx/tUmvQNeajuhqs8QdxdMsybrjBxBmeY+Q5YAc7j5ChDO1RxijhEmu3qB0myhg
FMZcMCRb8DkUH6/WWo236/dw+0SFUPmYxckSpp1uejTCnJ17lFtXXKbOHlHpTIiPliZdTe4OIiGf
bvJzgfTf507OuICYJu8XZLeNle/nyP/oH12K7xP+UrqFqS+K8k1PbYVGOr2VGu+Pkuc6Z6PIZTUq
5Q+K3GdPxqljPtQz3hVV0HtEHSgC4t+J/V11fKPTvfzRfy/n7ejDr6plupmRFg8JuVu+/nWCeSEK
5kwbUKYTDkN58zC24U7tbxcequoqTo4LALYi2lSStcARXX7ssRYDuo5+jqV7+9Fs5NhiDiaX0QBd
RonMGjTVa6ODCTCUZ2dJzbbiJpFLX7kNkX1WulrG26BcGVflDO0E55JwHHDfrBZjU1gCIOmfbTBP
+BQ3PZdG8iDuiEx2h5beSHQKer9c/wMwZtx2krY/Q/jDFI6zk/tXzMfVT0xfu5yGu2i29ShievQM
zeHlppmORfDazSYp/ndL0LSLoNtVgYqh4e/mRipDr7w6rRdptLaTetbiRJj7GGcP3BvX6eib0mDA
E+aif4AvfxjhErq0aOXIw2E/I/vlFhOH02GJ+iTGiSXMVYd3G70gmu0roLxJwSa83dWR+eHaMrqN
uzq4g69WCmvghZalcN+dv8WGo1ClgC3T45gtmCy3JgGHvdA9DEYxAObrj+dTVubzRz8NV/3Z2mkg
oal1BOuGFlbDbyFLB+tdEKS1pBlmP3bTb6Ii1XKbtBiTkZwRZsxeC5mYf/PMo6KtxPQ7yXCHjZD5
r683TUuUgKdLOUfxdrXBr12MdXjOjQSyl3rk94BSoEx/rM1ILfxU5N2cuWZxOEA7acP7t9I3viMg
M2u1FdEEFg0arHhJvlvLfnYt/7Mzj35C0rnngddVj/YPpiXpiS/9IB2VROSn8T0l/DW+9AowoMnP
MhBRB97O3IejdT5OpAsLiVcnicyQ75DdszNZ0NOoE2682L3N4nyHUDzXS80VnTvScpOZal8RNA0Y
JLwBHot3SfZHF3pOVg4pWlRHu9g4pTPe70BWZazhiVzHnFJY1YVJCjDyA13HQth4Jry/7NVM/1QR
AoqbDaLoWywYFZsN/sLxNUvBAYs+Jp01ASgm0H6kVQzTQp1b7UwcWcGvfZrIJFAm3DcQrBJkRFW5
Oecr6ScDSSj2JD2wqc5ahctzA95szJA0g+dMVsFu207tlrVP50M9MDqa/WZ8yO03z7fC2mJJ4Roq
As6LXJ9PRPmpzpivVbhh9lb27qo+CzPMbl/5vPZ49dIJYx4fz3C4uIAzFgSf3I60Y2M4aWeoaHH9
LkkCXa2FROeFk6Hv+LS2ZmbBcJsZYIqfNJZ6KYdlfjkbXi9gj3z7jh09L6azIAnM4+RBxbyUFxr3
ZJXXzRYhFgQ4uPuRbXbsB8F/4Bnc6cnGalvGE8QNYlnhptnU2QKsBOiEL7lr0I9emQUNkEdcQ5HB
ClOoyVzMfo/BRbDcyocNIPH6pD7DO0VVsNSqHPG7uGOHf+R+Q+dc3IhPpqoLT+fJjvSzl2dH/dP5
Lam3Niu8IvfDQ6AuvkohvK7PdnNdLezRkJxpceOSlEEcP8Nx8oNZAs/JZEl/gsK5I21Y8PlSuMhV
nENmy1jERrHsS3+frinfNmMwq/neSasL4iC6QhyPGLwGBj0/NKs1QBk/E+Xax4r0hspCfdKNnOe9
HkxA/OuvIG2MTzmg0+4naL2pxO8qFSrSHAHtTvc4V7Vxvh1Cxf5baKuumcHzccOUBixc5ilUOBdI
saUo154NxkLG3WAYeKPaRS8gl9VJlID4UfDkxI+Jynxnio2Ga5oqAj4hqIYKEx5aUZe08a+JFGun
ZAi+5IGR8IL7JGqCEKbemw/YlAF4hnIxgI0fbgchAdjxy9bJbQH9OUUZn5xHL2mPtMgaNr7vUr/8
A3AzTeu4iB6AW0v6q3IqKFlxWQKGbi8I5Nl5T6fRRLCrUbtyPPaPmqX+LeZcqRb7zdyMFq5wRmzr
wRG5LC7WImNeIq9ArxIoJ8oHnCA1JWBlG4X7DodvqjLSDJ2oD/epQk+NpXqgia4fwHKk1xK9LcjX
rMnU/Yan51JMcEXClCHEjsr6bnR3X51rMsn1II87GMnD6Uh3wsF8y6s7RzHsfsZRi/AMJQkmyu01
KJufg1Hozst3FpLzS9gWgFO/Ho59IhAJPz+HEI7KsoEPggsCIKj6IlTkWEG2vHvidD/msbH1Sjxx
sWzloCoemSP/JdhBDBIrmTPnihhi0uGvfVVDnIACVAbJL2ZtCAAI+i5A3iovMcYYzpcJ2tkGP7je
140eRN8taoU3VV0i1k9bps0wwXv54eBUMH0uOy6h7+JDLjK9tCf9+rsM/c7soKJpX+7uqc7qpqMk
m3RTGn0JtelsjamhSzn/A/2HHMvYS1WXtYg68i1Ruo8TAc6dgfy3LHejbtiqzINUd9zl/iRJC+j7
xFlWq5mzzAjsFrcMrclGf6EQW+tkRdX1cw37QjXbrP/cXK4QpDRUACk88P0x8dW0I9lJs6mp85ZN
Xbhvnibcog+xK6z8+XVatCdbqZ1aI/iXB4yN8HRCdveRBxBVyNL+46ldyVcYunPWxuleKLlrz6SB
lPxRIBci+TMwFTlKau6KTfTWgEsundgibfREvf805RV8c6bZ48pPgk0M4h2G2Ow54sYCeJKJpIHn
IaMx5pkAPCGav6Be6K3/U1eBewJpLEvvJoii6A4R0O4uChkEL7nsrj5sKYQj7GeL08G3kzUSyprV
LOsiF2J+KLWqyUkStS0NWd5i3PzOtWXJZWNZAmyB5SYqeZFGXigmxp38hP8YrvsZhbAuGZM3tDi9
dlxt6CELV8DxIJCP8vQGpT2PjmFh2jqe5LaB6jBBJv+w8eBAeF13iUwx+Q5+ssLiuE8Z9idn7nr0
kX9fLFQOOBIo3tmK3KPr9pongCzwgXH20Btex2HoHgac/MI2oxIwTUgHTgJKFtwnKyd1Ho55k/zj
zZUkrSRGRxMbEvtei3dHXyMMdeV5yLLXSv3aF3sRyGzY7uPlBE1IHgs5XDrSiicsUNtPIko/Fgnk
B0/aofa96BGPf1zQSB+YAJ9S98S+8FBnDmUecpq58m3Xmd3dv4wiFwuqmzwx7q3MQgIBJ9+uT1cX
Is/Lma/biO4hoxl2kEaIoR44QGkTSlWNzhVUCdVESqpGoEQ6D15E5nwpbODlpQSwP3z2T7n05Os9
Wg/2dCeBpLj10TkRneXUKDwvjuFW0OW9pF8x5HBXTZAC4yvI+nzyNvaSA+YVCYLuSJ4oCopIbNii
sP59hdr8KdZh3n8AQHu6MF9YLTdE63CsnCs6kZCqF4I/ISaqPHChVrZs3zH1H8JcTC6akBbdE8Zz
WdxI9GXPQsR1Uqqz+CqJphmu7rEoX+xOL5FtpAfzNas+RQS4K7toYD5+ijVyKDF37Kt810GtTJ2F
7JLRMXBAY4yNTezvwjeXCIGVEMSHC80xwcezmEhVrjwoeju9bkZDLEZ7zy3WBVQOKS7ws40Lz65J
myQc4JXgqLc2UA1FWb4l1XcC+kxuun7zpbAoPhO8u92g+cDlWDzzIV0KXIJvRNia3yl/Wpu1H+gc
187RQr/Nx7C1LJSk/zGnMDb3oIs2+5hQRiI7e3CpzIP+7VNjZvQxoAh6JDfVMcAwEF/T1QxhE/N+
9q6DIf1WV/mEcUoovnsprxzhMME4opr88XJuec1X2CD8QlhekFJPvzECmutL4EL7x0FWpDHlsyhY
UHKALMeeIlsh2kNODDePp4Zxy96mkV++MXKwiq2E+QwR1prSrI5boxKUfuFJjw3GnfI5rpQ6wwYO
wbHa9+E4i0ghe+hygLvYD+a3+JWpcdUvVPGR9C3HuGnaHY+f6MVUmEkCprFml0mel4oRxyjOgwTQ
1XeiFelhudvTbZ2AvA98rmLiQZYKEKkusnM9vWJYGo6+O7uyob9ZyLEm++yUCU7+SeGUOTQO4NYJ
rDOHosxJLWMt4SWZiLxBqyCxETJMnKm8ige6NNSji1j8DUttb85MksVQgFee6yuTpZZbfPulibgp
N5q4AsFo/OS7x1bQR+6bXhyGSDvYPnUqn52Yx1AkVASg2h9MpnUZyfEYJ4XNWa6CcHdZ7FgCSwz6
SLXjX/wFywTC6kJMqrr4MayiFQGBTSD0NQNnl0TGGOEAZ/MC73xAInO1q/urGOIPg+HYYQWSaayw
63QisczImS09+V8ZEAbtbMf0Vhi6o49hzsrvSH3BTs8uHynfNpy2hHeC0xEWKfWxT59RMSidDAjK
spVScpVZiE+u0NWYHbKRGtDO8Sx09gjcRta6jIlo4BCROwuL2a0pqsRkb11Wp3gAstbKK8tPV++O
zO4fRn1vQkVgsxRfUrgIUNmMuQHQKwETbAFb843Ton8LzNHSlqVywGxVfmoKhF+S2OTv877WioKG
6vaVFa3H2Hu5TZukHW5WsMzrbB/WBrVdW/P7rxy3Q5WBTCdcnoGmjtfsHuNZH+4zw9syNxrMlds4
FTylYXirtNu7L2qlgZVWK8SA/yKHpFtB5hPgJDNHSfd48FEaENkGe0GPBzOkbIXcIpgvrJ3LPOEq
mByDLwizQLKajuZWlXqn9MGL1fQZqbDMRzw+UyHvL6wVGNF4CugMz5seukt2bFI0h/LvQPxhjQnZ
l8ejTVYzuE4PUabzkrdC/+dOTs7qPDynnt3OG5N49GSxH+MTO1Jrt4SIwNWEJtVN+4mugqdQvAGB
qTxlcpoaB9cLwxX6EOmNo4lRHrWRm4r96UDyf+p/bm5whtdy9Le056Uec9XR0KJfOr0RROFNkJtm
d0F10+3vQFDjcmMAO2WdZWlsmlF6ZJJhuYoR1ntove+nH8XzZjbg5OSJqkIeXxgvu+Wr/+QA07Fb
6gcsUK+8r2zpA1emEbWlHwA6GR8Mv/6Y7+VPWgtvVj2qdeXymQc/xFmLBD6OPRGJiEhpSIWo8tzD
QrTJt8y9n7uf6tCLS9Kgb7OdnZ+RwK1exYiHgYawqvZNUhV0xliDgIONFwVP/K1C/P0zFIaq2ag/
su/c92JH/VnfWenILB/YMibgSPjY1PhbwFFWvSUE0eEcaw3RAS73owJGmnPVOK0rV2783R0ZdyNW
blXXirtxk0JTRU7ZQniXBKiL/hK4AwghjMaO3rQSHvas5s++C6ODwrNmIA6LQAUqIUrsou/b7jdt
YYm8zkxtWL2/eeJqpV4hs1bt4T4xl8CubpM6oQGeaq+G5VvD/D2k2olIfkJbrKvKE7+BAgBn9cao
RJp4zYMt7imYJmWiGfnTbHZP1uoWMriWEtU0jWa9n1RW7+fNArkNGVh5sleczlmLOFA18jgE7Ukd
d89xZU0MUap6wKdBjLcaTIbItNBppJQDCZn9Z2To+dfHmRrAqabQpQSXxsK/gyLdtfiYS6apcqfs
x26wR4emsRqbdU3o7Bpt9XC3N+rKYoRpUvdX8zVCXQSdXHH6HPcFuOfKVqoM5XptvIdDTYbm5tvG
yHtZydAMfLSXi+mYu0Da7U3kSyDUNwbmRPuUhUI+09VmFJMs4b60vazHdFLuscLL/JaN0kmKoMM8
RTTel7MUrg3PzeWbsCxS32ylmLlpqzfLftGdOzcSaF2IjngwMTr+yLL2i0o9v5UBj06W4SVs1Vea
BEcqPKcf8qipZ2nLtLN1LTq1UAOZIoCrkEVVGRdUJl4AFzrnEIr9jVShOBjn5hkofQopuaBbULwp
iJMRULiQVxPQMEQkThPEzqrWgANbIFP7PtaWkSIp/Rw83fGiwbxTO+kMlUHwMqPmIjn33tJeYGP9
3hKYejZsg76euzgs4yumSU0XI9f0LPJHFO7AtsxEkuOhQEXiBQgWxqCCw9wpopX1SnzJy2vGbjRJ
SHJ1CzppYhzyaeTWHKipVVi+TImAXMdO4ZsL7T2VfjICT8XUj92z6ii5nyGBCgU8CtBfLteqbDJK
Ly+tEKNQHX0cfNOHFxj3hrBBKpKty0mab8BJrEdeUwyWpovh5BiDfoGjkbcKUYYHMylI28Q6KZGm
NcQAzeYMBG+AfjhORhfbDnzoEIZ0ykNfJSvLKfYg+RMDioqL6uUpia49WoWu05jIQx5DHwsuRsgR
Z5GA63TuHOcdEddsvWS+8R7yhGuT6KDeJfZqs/YBy+wJ6FNRPJFM/pmz9JpcLWTvm3UcH0rHNCLi
AD2dHHTuxioQm35cuL1fDA/uXG0sHCn+Nx9hcBtGTjgn+p5gA4cUTU9hz49SNdXVmaAQMeqTi6jW
NyRlrlClarZvxWoSTvFGq6hmk0jfy9YuIyoP4V0kb5pNQDkKRg8e/Th0B4st5M37BoMK2VWLGcVA
yuWLs8X3+2jjS3tbvzu/vTjkhNQH8g2rDUeulGH+qOQmktT/tn+9M+3GuX0ibbRowuF3z21ESyWG
MQt9h/wIvkVzE/9a/tdMVP/v6GTccM+NcJyWmsGudoxDBwi08kTeNn873exwENqHUYC7WWwmvWh2
Hfh2hkW7DdOIHnVYe5vyy+Lco0KSOzUXd/kHIElT6aWMlB7K/m+ZJBBjxnhY9EquzIwTvdr73lST
jaXngwQQ3A7BkNpSqFJqqeByXZrK3ts5wbaZv4WGwVlL6YXXHumn/TnDWrbGpe+yRIUGkc5CuAkj
5f2XzTN44nxSzeh/MvIvbxiSxVky2O8QXsiz3cC+32K6IzpYL0tQF1AD6RtJhRK8XVJU+VDqq7Sg
q5zKb4LjMDrdzskVbE8pqAlEFsjO9D10GdG4TANPWXdD1LHFkwUgqPQ6Hs3w+0FxdmYYpdQy1mZQ
BQ98Nz0PASOqmIIwWrsZ/dE09KCKvWhaCjFanjpZDo4wmNXTiA6icbkXxQLLYdwE/XY6h4Dianze
jKYFAEmtzChaL6vkNPSMsuM7HV/t0phXXz7E1v2IdeOKY1nUjMZpMlhbrG8cFbR59ld/4sJPY+jK
kH4aftcodC5TlK/EPrncf5MHj3m+kiCPW9pes6/DK0n0S3EQ1WKBOkJ+LlF6KvMiZ5uc4Ppf05NK
Hgia8W39rRu6n2zn3GwQi3oVg1Ew21cr5q9IkglYqaaDvietplzIXEAyqUPWubnYUOvi/e7ez1lW
CvBZStEtP1wtxjKV7J7/V/6QPkscXT8d4f9Y4ao/leqGgNKRh+9Ovoc6JtZoZm7qvIl+FhOPVXPt
yoxRzwQLqdT2bebqP1aOnkt833cnS5jN67bwVV2iNIMbFynDRvZJZxLH/QWOng9XwiqbcdAbD+A8
EEXopoe+nx2gLL1aWU3mHNdNEjdgOxah7xYqmfwcakdncmhFuX9WhJbnwDhENEOZ2TSGaO8EINfK
rlVikHImfj+CrZQbNUi6Wfpl9t6/FW3i5htTCgFA7r0lokMVyF3FgAnofn/JepMCCDdtngHmPVNQ
BEDNCoQ5twEuHbNyudRgXg+arY+8KINuV/jtX/q4oxpi21c7SG52JR167ovmEheoz65ptO702mQO
KJBn2X4f/7jRTLPcdSA4ZegcnkPBKwQklCGD5FT3rXIBcM2lFi8tXIAJdzZof0UVWAmjwtGjQy4c
HwJXOAKCa52g9+OjXQiwpQLY/pcJ1EBBooWwfxZw+e7fXmcngvoeuGr7QZlbVWBUG/LjnYemjZVe
9Y8SkN4Ia2vbI+9UgKN06x+5lMEa4101MFoYxBk8z0mKTWXN9ujHEfSbCNDprA3N5a0IEEgNw7wI
BXQ2XgpmvB8IeOHDecQ2HO6yDLiZnpISPRsBAoJfkzfk1FP65vTSASfVexAvfr+1kd4hj/+wKIOu
wgZAEjRxZhChRcxQMVbL5lOxK83MnMw03zhQQGfWqAkOgxrYdu4cjV4XPapqlj6K5g8SQIXXMdyd
iVEHVgA/bBgbzAvTCiMmFpqZh28GkG7nsQLVRy7yZIay6Sieqb4RBmo4gmULaKBz5lF4b8rF8RWi
Sn3IcfawBoOEwv80kA5k7L34JG15GEX3yI+4bbjcFjrNQ9Wbfqji0sQtTPixshZ1MjftYb5+pFzZ
ZtQIWb1IwqnTQvpmDn3/o118n+g9xTa/+e6PyYc5/Uher3PGut6y/xfQcF34fHZRXWvvedHhVdA3
SQD9Wz66Pn0q8taOa6YqHdLMDKhHJ25+puL/zALsEKxlwUuXOJ7kbJbiojFssqnaWPyNrnUKRuOF
XI/6SB8rxCKoUy1j3CWAqFyv3MlDPkz+KGxhz6/N8OCfxfa+CRlkofts6aABJlqSG8MRJEJWqz6S
f3RE0+vSh+J5MwNhspTdiYEz1MqYZ4YYMPk8BWTvOU24rGBHxJxRyg3sOdGXwjDGsHg8murs9w2z
2rtT5Fl5nvmZvlUNJh/j3vvTXnnGBn9T44svKkz+X0qLrdJRwDawjbSlTbAmMlfKtuJHnu5yGaOg
yipPjkDQEPQgr8q3H+NHKcD1A0gtW4yD7CBhAyVyJM22ena0aBkuwMbDikXM/SNPPDeXlG9rhIv6
XHIe1gLZyOtmURpdyHuJwiHU+/vn5xj/7pWTyt9MHzuFRb+RMPcvtyDj3jQlcp2iG0Hhsfulnc8T
rvcBmMT3jn58qN1oeFmhjL5CzDoO71CTACyxxn/VNkT+4N5yA32D/DrLjYU8fqmC1jgrcWvw/BCc
rb52vabaNHHUr4OqURJwI5MLia3bt8C+GBPvIiUtTjjX0dQsi7xnKF7AAa9BPZC2B3jAjMXmxPPs
7c5Xr1U5ESY4WT/Wpt00vtAocIHsuVHObpmU06GPFm02iuJNRmjYIeNhba9Th0zvTjwQz7EBInWW
aswGP43drSMcZcqN3bC+h/EE8M+3bdlwg/vqEPekja9wDaydxX9qSyQX/2ayKg3NeZ0FmbkMzxGv
MXGUTBQiiKjC9+D1IplrV1nPVxTJTspJPMxM2GS1o4cVy79pU4Xh4uVZI5ik5dIanOuDBAdE/xic
g0orp4ZnNi0rLsm5JNka2/+M0GOWM9dK5qn7dD2exhaeLmbEakauleT0VsSybsxuJarCcThnzn0h
fCQVzQfcW9gIzssd5hgsdz7FfkD0ip4M1fNFHSZbWDvmAsk5wud/2Z4BOtEyzSKsvQD0TtXAqA82
TonwIAISe0XwareDZAdShI2sOlTc7vZprjwc0jfTQBeL2sp/cFCZzatAkwSFGJfm37EThyzH4cYp
yLsdTlyitcKHfrtf5xEPhDdM+jzKru0IXugbjVjS+a51QJZhTDfaQnFPhz5pZ8HREphrZY7dvdGR
/gl/8cSv7dbetkw+biwC94OBQBZ9CRoJrGNE0LTFJSZgQBUnRewUK18208w2IKwmAjwxEu6bocQI
Db+pqimKDy6pSkVBOR4zPrDR1buV/m28csWbOoayy/PJw3Kc34CwNm9crHUZkmqoSlpmHa8Bcp9c
n0um8YA+HVERcAcYtiluxKQ3N6aZiobdM81i6l91RJAJ7GSufXgYb3SAn4oZWKEpDX2UpEJ/uYi4
dbN8nQhsljw7AYFzMLV18yKZDootgXKgwH+OWQyVPk/tm6ffNu/M1ZLYnM/+Z5UiiZIijL22bUy0
DnzKn+Xv7aFRWKVcdOdptnfsmq3oiF5AI2F7tSERfsADwfXA3ZmGUrDKQBvb0XcCYScek3fxnjXq
W8oY2bH/IJSNbV4Efw/GqjD1omUoHAbajZRu0JEMwG/dafgTFUFK9c1XSbklYLu7h1VWvVFzs2fh
aMHayUKlj01TOx62Tj/wuITGvzJuRNNkanuyuT3UDlwmPkGkbs4GdMuly6n840ngL2EMdk5ZQGpW
eNVdpmzdy3w7+9T3DfYN48BYcOt6+EQ4HGjluLyiVn8GI2ayYv26SKTie3woFgfCTDpdlUcxJmGX
jUVab3klhe3ewsaD0ZNiMiNWYt6ODGFrdRxiz6lM+B5b34cnzwM3KwmBmFKOi3SASeqYd5XVNiV9
K0LMlwMWJVibyg1ZaZO1+6Te4hxK7yiQeXDrHYcJ4kLl9xf30tomYlorAR7F5bjQd066PJfaX57f
k36cVrelYkV0B/qHM6YA4LOwvA7dNgG61c20IrXwF26I9g5xfKkx9M+UPfJDW+hXG3tDitwUrRAw
uI8lx2maOtYL+ZPcTFlUTrdYzZA040qtdfZDPpC+0Y/+hL8OQDumpQusw38Ia+/EiCnxSmhW23cm
ivBZDw8PfbL9odFTkl/sao0ycTo38ERe3kfQYvX+s0JG6zkEaX9fnBDsBf9QB6AmSBglnl96x2CS
gsxMty7DVC8MPtfneB8/Bsbfloq3Q+cu9UkQ04Nu7KmWZkkfVhc9zs10lv8e5YqNWZ8nnlvMVTPq
bLqR3z/zsLkYOp/iAILbUWn6v9OXPyTemkTiTG/zkCgpOCJG1q0YRX2IBCm/M+KdfmU3xHhOVjPJ
TQ0tzX+PhroUthMuAHNifQiM2SbIL8aMYrbIuoVMPOSWOhu5Z1w6UFvcO0p/NWPkdHO1Eh0+DXzO
kjbyEjWsG7dcnyEoWrfpDXjwC4iOsP2AQPR1dc1fLnxB5nvSx3WrQJ5nmR0IoIBzl6uvUjw84bca
HZNKz47UkZQialjTzIs6R4u+5s4IZVl75kmZOsqrnR7q7fqAvBw/G3E7lI6/SlZ8BEZB3PiiuEbD
OAARlUrcOQc4g7PcKVcUYnp5zhaGgHTVGDKi8KmMy4a03I9e54Npbo2Tjtyf1Y1mrL7vxVPJfPEq
UH+ZRvTa24jmWjNk3xYdGSb995J6VQNFdAP2u3gj184PQQ78MTEmsec2Ihp2O0xwXgcleJ+j5Unw
q1OKnVb6B7SH+YfMf8hdPMjewrXsNZoHMArhuKpyWG8d9tvwjIdSADJ5OFgqkjqYMpxTVeXWTYoo
lflwHUwdf6Kcw2k9gvsIdBYuO9Z9/85xzm0nPqHT7P97rvY4vUMAfADIjfHTFTZqaQcv102Uv7gq
6G26wV0YTdl4XQqrWOqqXt2vhXTkYQQ8G9XMg4h3JWvmdGAeW7XoX5YopMO7LJm2rNTnXkxb4msT
eC3qKBpbOeWwrdZY1TKqgxRkpzvGZiZzwFi+X9XOx2T8kE4NPl63A8iaOV6BxK/ShtjnKnjv0BXI
j6wOpQaZz1LzfnJaI8C8+SwcE3VxdRmOD3vpWhYypACrZZGXt4vPdDqnKc2mklnevyPzRiZTs3g1
Xf7WEUAh3qGWNkMy9aA96YMVbgCRdaRff7w7LyCTUFEBH5RjmajCt7U1JfsXgsfqkfRcZgemeMjS
n8n8HSlmTvHayyw8pcRdAWAVwfGPxhBqD+Sn9KNwug2fULEIgYL7DhZIgz1zAF0Xu6uBsniDjzG6
S8IsU7o9OEKXJEHI9tOMalvZlTSMJlbvsa5mbPy+82IGmIjCx0U42hxLS2fhAeVrd0XKqfyIEweL
ShR4bd0VZI3X5FoMu21+Rs/yKBZj9RhbvLN12+u1T7CCBWZOto9gDzJ6wO+ouEZ2Sl33BSkT1fJj
Zd10HBLMUWUCxUjrc8Kq2LAdbkFea6JVD4uNJFEl3hueCNPkHBMVJTd6LFqma0Z6BakOoUwX3gfX
VlSUZILzFHdfBQYYr8oSJuCoI4FHH10qIr7TZJN5MX5AiekoTa5gDL13+6Qa28W5mJepUtFhA8kW
xToVgQGu8KgltfxnVemgf2EpRe1/nR+SQpt6rZDBiMUMEqbZT7XdF84TX1x+6W+2TxBNMxzO3AAH
sEfORpJaVxIyurWCwzVuZritxRFlSJjQAW2ijCFej26spg+7xPEfxC8JBb+zbOLLij7VuHD6o3yH
z11IiytXB9di+DnCWztO+toqvCj20OEBNmDQQrwEaLHTF1mAB6/5nwyJNqToOC4o/1+WounM0Ssr
nyJ2CKZ//byaY/+Tzx4I3YkoAVBffxut9TARmW06t7/v+BX6VRpQphBgBDaEgy1BWJ6IA0kUlbeu
AzEOdcQuQng/oLaSUHEBTpa8d4twgfT/Cz+51lyXhVqs61R1tZNHK/t/miWiRxaOTtceQIVr12bg
0dkBOgwhEEjS4ILYuVg6Is3dYSPNM9iL3ORFkMRxb9chw5ZhjzzTVUWUAEkmHa4dwSe0gC+CPhef
9jvi0Vr27MAzTBKX7rEJKDIYsNr/uk76SWf7aEthOuSP3KPTvYke9j8HZcxtBap4LAfvGkZ/ftq7
bPq2Eg4Ev95mV2wrLvKCJxdEQErAO7cMuImrHd5CFaFs9075HvXT3f6jwJfEDuwXGeZac8ExR/El
BRnPQUbFT8yQVViQrYGjsHYnakLYNWFUqG1iUR0UtffTS11U584y0qLRFExK6f/68iSH0jMqj/tz
R1cX81Km3TaV3NwxElcecLBh6rW2PBs4ziSz9hiGIrYw6vdPiasZ3LY0NSucgvr990sKaXmPZGn8
Xc9ikoK7SzdeWGrcyK2Kbvx/4m0wSZKhH/y1PuNdZGOX/i1Wrrp2C/ouWWqtfKqQLfYM20Wivc++
Eu02ahIkkiFJWQyrk3QLC10PHd2E3Y0QPYoBlyEVm45txEyVqCLQ2UKS2TUM7utH9l/9FvmaKFqP
GTy0V+2zIFdqqVF+r2zCbB4vIdyy4hAyQRBEOzMvTzTOZMSxfPzuhNkw8v5myzaBsEHmd5reNcqf
eSdK52LyG25bMUSi0njJ7OQaVE6Jg/KSTbRKwJPXVglsB4Bi/MZBioOqIlDKVXbQcpKdMZZ/z/e+
wNAYRatzCj6WbIEDpqVOC7CKjPX5H547UL/qeMKwCnokCB61zTSbtoU7fpUnUhXy000LtEJdyMn4
H41RiuOrynO8+7s9pUYD3bvQ+HRG9/0Ny6sTOoRAD8RfqW2Y6L54+mbcNzgXPi+lC3vqxapX07OT
hwIDnIDJSRaMw5n5nB7YZ59o663yqCYUkOjiSBRDEF3pTKLO/cRPHGIQMZsEfxope12ChtrtRzh2
IlYrvxogLmlH8+B3rrLFxbrYJO6D17SMzud9Kd57i7nPqZi5a2nirSnhyFWBlFNSCd0YLDlR9puz
/eaThPHRfaM0ZXWBDy/YF0MA3YbgO4K0jKmsGGmHLdeNDWLcSQ8jTxR91MFC6H1B8SGRk3OXJ9jJ
KJoqKczUU1iqLk/efRVRJAYmRpPheXfy4r0fXER38JNpQI9VyZ4HkNu4wxtTj3rMNZujViecafdl
5QBodemwHP5Ra71jSo+OhCHGgPZ15J494Ck8xpe4Hs1iSdij9qxDRd/2iKqGITRyBJZoyz2/isFo
YKb6mfW6qaVP7O+uXEG2vmOz2fDNYwpNIUiy0Q3ia4zOuMSxYBvYfhOks/MnJzq1RtJQaj1VV+uh
g9Vpcg+Br64XY1pjdnR9Yr4aStJRmuyzaDzdi2oGzH4mYRxVKEYMPtucPcX0p3YMEOBwb6Dn+1pH
AgYG2NfpcCeytTFjxQZgbHZ1zmNKW05G++248Var3GNLINXD87OBAqVNRIRttjkMmqZ3+nj8JzXe
XDZU/2liR4NgMt23vl9iG11yWV2Xdsfi1YqtU+Hy8rrgR4TZ6ZX9Ad3PO3RjFqMaR9HL9NSv/i+s
uAMUFCb7HVfTT2u2NRLBReerRSLptgSHbYL2Ib6dz5y4WOcLe4bgZpXj2i9YN/AhBShE+Jy04fc5
vZoYFAheJcFjD40kyIJfXaJwWb+V3NtexbqWcTS9Rf7GKi+mNYHIgbv8DbPW5RkIBI3+Ays2v1Dq
Yd1Fuq30X5AuvjLY6B/y14YLjbax8P+NA3r8fWcVB+6JosMoSFm/e98WHFTUPdgffs8uO9hwvkfl
N9wawjrPG5h6SBPldNRV98CeSr2gBtsENvyC/Qy8JjEmUVgQu9b+I+p40HQ/cc5p9RPduI5YjjH1
i3LQIq/SV11+j9S5DiuRgEakuSjoN9zqC5mbypj/9g7l72sIhPlNq0RDfnCBcTle8xMZxfk0rcH9
HpOhp3f5+pEcs2y1X+MOVHZ9hgRPmKwZzGxy5+TKxVSV9f9Rsi8VDMX2QTPWZtFn4X8Jssua8umT
Phm15xssSP+XZF/qFXg5HZhO9FkVr5VFlkdkn/01HysxkyU2qyJ5xSYFKwGaSOX0tWnq1FCGbvWc
P8Qy8C0Opg4tkj7nY2DArMhK3qmbLuQToCrjgeq1aH1lLOBxhwI6NyKvX9v4HgYA7ZZYcnT4Wb1O
Vi7Gp4ODjxlatc+UVnFspzL4lRfatWPVvFz0hR+pf3SQKml3+IFKhn3Vn2BHgQ+IJh2++C9OcU6i
dM5uRnS2Gr47OHjQv476ENbnQ82J/dU+92MxzQWnTVAQeZkNJxMiNP//S3v6jpFWH/kB0YHuQn0D
3Za5v9swKI0ZfLco7Dy/Hrjqv07wUKduJPDboXFsxLClL4lZZJsCuLE8sOoq89JBJ/xlJz/eO3br
h5vNvHB8NObUFNaE90lCLDIm0wjEyETs3z74gnY7UJ4Foqa+cXefPJMpdHgC5rD1dO6eL7PFD1mD
+p1MMcOD5ThSiKbFkIsuRmu/UWd1nchHV8rxQSCZxE8HTSBZNQqX79G+DUkawuv7/iGfbSKTPlA5
4S05hxol/bgluGRpvDm0YudHudnp6ownhwXLY9OYBruI7VhKa8dZNfnHCrAzYZKl+/lLwbn/fRj9
q3N+UUX54eTUfon4VAxtpQpxxBH/B9M2yX7jIBELE8yGXKRDEvDZi0zjN/KLUsdOD9mD/T+/SWUu
/QW0H6ApQiSCN82Cz673kbLN6/78a7CsOjRqtb6NWdVqGxtwYNgt32uoSj84i6CbwqwNEmVSTdOS
SG7wtK3QZQczQ4DCKRjFMYlpsOHYaoiUrzqVb9DxxsWMl2KgNzWbQOgXaW0RmO7iMhimgUB84gvp
Ysb4QFTEZmmWQo6ApyxKyqTygdDj1LTgrjgLzKJdeWp++zRy/hAs0DjkPiC4tS4a6/DlfNeXaWKQ
ELsmxnE8iiZmjcBauRSdqlvpK6w9Xz7dJ71iZ/YgSWGaUHfZsdeHDO9mTxNQ7WhQDc4YTJSSASz5
WPFHpf7HYoNVegAog6n0e2BfG4M+QBhW2DIbFZSEdMUjJmeD47ZDAkN1yKi3OOMR1Z17IGUHMr7O
bMLlQ5Wek0jrnlcHXIm1p+fVcAY3LFc4qUshwgpCgpMIiVfuBl9Ypqemda86GWXbMjw7nP5Ke2nR
o06S1z7+0H6F6Dv5adLT8MO5lvlQe+gHd/dX/8CweqBIDp50WgyT2oAc9QuYo+Lx6YdP9+xQxc3f
pwMqB4yFR+ylRpf3+eHA3TR7fhlk4yQ4OsvHcbGZQGI5enVUyMMpHqIDFWfQBWHVX5Qhjz/ZY6/I
TiWdybSd06qPaaZV4l0OzB+uNSd5P9Y3nr1edgTU1dOrOsNgwAJG0yRSP0gxNiS8HsFXCTvJ3X0D
/HYVryGt4KBifgh0WOE7tDCKu9nEr/OU9JohvR0/zaFDBhEH5rGF6c8/k4Zj5I3XIyPouMg9F+is
bguhCWvqdhJL1AhwdOJUAlpqTlIHAoa6cvIEHaN9NBFazgUHTrzlzZy3FwJ3vP7hAx6BGmeJAHLG
lp2HdtprLs5H0fSItzIWjvSxuMySCfywvBFY8mIekh5Gkk0ThtZLTRjWU10rreUaQMPIPwFKcXUD
7GOxeheuwg33AXWmmCAAyAEM3jJJ8xcdzlgVdZBR1myUEOiIhXgMBTNKkRMoKgfDgDqfOkn+Gh/U
iAnZ3AaLBUtZ8BHRJHCyaVB5Do687aEEVmuUf2/UPJe7hk/SXRhFss3i5wGWsHT6ORbnmnpgVGU8
NZ+XrLPyPZXVnByyry2nhpR0smUc0ctglqCB1ERTNijtGqQXelib1+btvQNUuqQrvSK/wyCCL1va
gZ1O/irwPbt6LlN+kRdYfcNGWjnzpr3e7z3NoWR3dSYbiQKQUtrtIEvjoOm8uO6DmtuASO54lmZd
J/Uy0Acbn85DK0RXwgJ7abIv40YA/VWin9YLF1i2MCUz0BzUDb80hb6NpmdfWBpVEtsnuNkM4/J4
QP+tnGCezgK3ci155oJ0xqKhO2yVG1URtFTTix1jfHtpnBzhE9OGawyiuxurpPfrlDiWuv+NmqZY
cVsgyA/LhdfGT4uazG/1l2LuOuzhXliSRLKwQCK8bCkMQRzTUz2mPega4xz/POUEYElw8PDdQTqQ
QyI/9ljSYbobBPHOUL3QaD4AH5QFdrC0Q08u/Qz/C7fd3dgZQwXLnz7KfHQ3yZa6LUrDmipu1SGG
M8HCdkXpls/ftzBOd4wv1aKqHY+sBBMs2EQ6bZvs5MKWt+JK5cFlvLO5sZ9YB9x73U1D72PKxw/Q
ZWX94zf671S2xnBvdxGkriwQ6IKoW6hWQbEhcZWCEyRzDO5lnCDkMl6NqvUw0gs5GbaC9qNJZVrg
4Ag5f3+VSxuSlahV9lEtuzg4v8zbgY+LZ6uDnj/lO1k1pEGlaPoz6W4E+oQmfbq/kMbNd9Baeo5D
h+IWpE69kIoIL6BidpstvRj+I/dvnX8bfOm99Ewvskaz2Uo2Fp3XZbwfe+zXRjxXC2+p397+REMo
dchQMgiV9ehNN9Akm1AP0WaO32vySnuNhapy22pB+tuMLQvC+8tJjqyB4t3rpxJnd44hKEj95ken
z4bawnX8G7wjmNu3dbivhpZ1yBFHM8YKNatS48xVSeKXiDwYWX9eDZDn7vpucHZB0NYdq3ST2Lqh
65oDrz2+F2MHhq/idxP19N5MomI84mzUdGWXvuuYzznzwtyw171hqvdwFyIUtPPnHAULw9vy0+bw
wBTinN5X8IdfU3PyvfinDeJAaklhKju5nqZ4ogH3FalVp/F0Evm/IBmhTsxLZhtO2VR2vkR+ZhCJ
7dhYD8OKF95fUVndZ6wuxePPN9F0o2i6W49QHnn+qinSrl7h4+SMAyTqAgA9fTYM6R2MVtmD/EXS
A8doNgaVqbSmsHUDQZjD9EY6B6HnLifEioMPDlPL8CGXyH+/mZIUOD9jq9C7VHYWirgN0C6BnjZL
iekKkS+qwTBfuvRR/9CKE00SCG9mSXQR5pvHXrcJIPebcLHEzAA38hq9CxbIkOwUjIaJfevIJLMO
xai++O12S+bfyppUdkyFUqb/ZSsI5EBwwg3iIo4nhlpLRsa6GpoFfA2CW/Q5apQ5vIY6hH47plB/
X9VfIIRBRy8ellA6YgaFdZpO3afWCnt42O1mQgjIaUzteAvQctDZRLZx+8y6lqpBPU3s4YX2R5WG
gowdG2/2AsiuzBoMnqdCHLYt+uy0rW0MHj58I7OCPEW3GN64ZwLbf217n0hffxdvp7CswJ9AQ60V
hTcz8q4pp1IBWeEqyKt91PWclvwjsWNQKpwceC27emlOsGIuLzeEeWorcz1ObNM5oRpt4o0P7ouQ
pKYLn6Rncfz1ZIvYJ1T0gu5ZUgrWWGGzU8PIWf0766l7JAm7hQKEEV9YWIGCbc8K4iBqkKY3eHKM
+2Nhe3G8htW1P6cwHZyAmCpi+vAwL7v6gTpBc2v9k41rReyYOf4D1RnrgWgaj9LoCAiHFNlU/6Ju
qa4Uq/qm9n5Nx0yEmGqHPNoZwQZuuzKTaSiK3PskGs/9I/ErYyn1CqKcHq/h/bpa6j4MpI5BpzpR
6KflZBS74+tQ4Sm64gWR+Jt910oSyaf8516ZRp7ejmD8ugdxB6WHXljG0wvjxEBRVjOhSJPW5at8
ANqM1Se6TZY3tNx5idw/9GgyRBzpyB2GZOh02pLN33/Zo3o9fsUl3SThwUSYvaklxv6YIv7DxcBB
Qig45hVWICg2LS1ZD4sdtuqzSKV98zCE3e/JQJEgK99EBVLVXGnTagVeyCelW2ac5VlcsITD6nJg
auNhYbpzUpMFDUVD2fTNjCYKRqja6/wD2ahI7r/HjZC/L6WIUv7sKIGNK3YfoFS7vbCKwRQBJUJB
OXPKYIq1IA7+DkARY/cOBXGZ51hwbgZPY4f3LVQzrsX1J82g7ZIUp2bGu+V36Ae5cCrNkWJkPKDz
3E0wQaUyJFSTrmP9Sxqw9qQCUB714+O8qCPRVRRXE54jy0+hctog4iUl61IjjtwbO0HGZH+r55w1
vz3pNIFDjE5Q8jnH4o9iTOSjt6t3gBR8iX89XsWGtUhRpvFID9XtzMpc8a2sRpEbXxTNPNp+zEGx
poSqq6tq9UoqZ3MECXwxb5nBnzjGOYSpA7y8OZQOi+0lZgKoO39BT7mQLX7q8VZQcedMiJIqHWr8
/3omMplCbXIrleRpffYlLJeJwYS97/0ZCiOEaewH6UQBPircn4OSxvL1JLn1/rUQferuI6dSKa0z
V0txzbB4AqhI3t3i9lIGoxLIIlUxJoDoVOBr+qCj/OzfCASYlymEtGhHhRv2oeusTJ8s8MyyMDkC
DvLzKHfLwFwrnAeVBJf2cB1FUTce0XurUI5YeEB6fdb7n7ZQFVI33uiNUyQBg7Oe9V6rzZ2lojqw
hPglnS5yW1UOZk05ecEAF13pWQhdLLPM+ESSLnD6FvFRQVIcM9dO7RapimYl1iAFwsrVVDepjzte
Qef1fyV93dZrj3lIV5bS6gI+UfT5q8PVz/Sao0eNi/P8EQ34jj6vj+0ZXgICirj/25Abm5jjjG6k
zRnvQ2aP9fv4SCtgwjFBCY3PeJB+3igEyOV9wMamy4moVmjaN9YjmV64dqkhkqHQenHx8pFi9N7N
lK/cvC46GQTi3Q/7IU5KdmyZXBQyJH+ot6qTRtZS49XD6J4BZ2+oL7cyRjsy9ndPkhNm5DtvtjTY
/PLZF+8t9WonvvxiG7Hbfj+tLfJs3Amixn9RvV6QtsGqFMatml8y3Q4hZ1FcrmPpahUb96BLfziP
YSXjacOO8sABR1DWLikOGjNOBZwaZPWIra0JoFPtWVdl9WqBaqcNsTnZ3BI2pvkbtPWVLHxHI/GV
+6BeHark27hXUfj25oZyNskDnDKB4DuClLofaPB7gcEHvTO0pLpunxRyviGKHdO6xb/puMo/0iLb
WD3jI0MbM1+7FcT5uc1CrA74mquhbdOOX6gJIhpCP/czluJ64hGDfmMQrBC9tDorryV7N/r6ora6
nu2+GsK1N261xUkfMXIRO6q6cKow+BVCQvlSMZ9gEa8yjG5LlROb00W14phIzxMzPdECNFnCtUeP
rM6WCyeSNpANcvs2I9LFvxfTSW03rSwMrRW2bqVbiBqXLElzcxjxT6WCEYaJhpOCXJxC259RXW+Q
NhK4C8UvJoRri5QWBRTu9opVUa8MU/nWehrGSPK0TDeCJaddP8untf/jxXGumYQLt7JG+swGpGVk
AgimT9KCZW/UsZdiTTqmhMe8CdZ8wDd5aGAa81mYFPU0pFaxR5s4DHjz2SaaSSGbfeNmGB33IDKW
0EQVZN1G39MaJSMl2J/RiOYSuNHZls0fsQmJHKTrDUXI5APFSF7b79EAD5lpbVjKNjPYaDk57pL9
GnLBgLw3kEHNkiawrN9TwU7iJZz4+yXL7PH3uMpAIzUzRQJROXpzbHegxZrC+NxvDMEmC2KTrNwe
oXqdDB4kqBvnH/VKJEai0KyF86bSUUV1fDfHdbvcCZJKnbRue8KGR2da2u/x3ErVMRsiWkSnZ5Xp
eLwifmH6MP78Wfwd3uccwwGiUJdRsjaNMzj3RcI1MqMZEwVbCU8y+IeLdxu91Mrijns0PCj9mBQ5
mhprptWL8DB+HvxBx7O+pc0o6TRNIVYHRh1ybUfXJGbJumgMiDfRr3yNuR381Rag/2JhTwcaYn69
exxKiex+bpt3gGt26Hd6NuoNC0205vNXM+d3FnNUv4Y8qFjmYwvIDuOOxhdMhZa0eRZUaPIqaMT0
kPnxF58LD6OSbdIw70GXuhtG5z7MMwEJqiC03FuB2ryK30PfDe4KfA7OCwD5MvPyfrGYxdyukgtW
xVoSz0fOsLeyCKa2TrongdVGmjHhqaKHaD5umM06rTyDU+NvhrEZ9QfAxVOUIvqdFqH58pEzJpTT
mP9YMs2l5ft9vqFtiqx+gD4UNO8Wl9GPiuGjmpkzJVE19CKFPngvol7JHMuiXfsw0bntCjFDAwZp
o9zKOjG/dbbvXoaI30JR86h3wNFG2xGhRMI2o7gVEH2Lc1OXHEoWeN6GofJIykG7+ynXFEO4B4kC
9p67vG5gE8Qx5Q9ukhspl66CHbBqAquDPwlx1tfRvJybABzVjf0+Jwysxwut5IInTDlRob9UhqAj
BDNlL5bwvLTBO87ZZlYZmBBLbOXk4+0bX0M9FjT1L1zrvIg+5t2ipnoqGTsC1C4q44E5I5bIcXLj
64j91qjB0SY1sJFvI2qjVXQ2q8N1RmzWgPnpaGkB6DZ5vOep+5o0qlS9kBXtnSOx6rqdDK2lwLnZ
7OpmeK+BCL2evrVsesYWbKPW52y74qMBw5uGh5SsT5J0FVCPp3ZxlmVSeKdEEqu35Bk6lbO/Hewa
qLuG9vnJnut7SO8W+2TO/b0yUxXzq79W0t001iZKmZcXH+SV41Uc0OcCcASeQjMKQmSab1+1w2AT
2a3PVQhDOzslaUU3oDIV/W2dE7rvDD+gNZ1LCRnzr4Vc/wp0m8ZkwynhOW7a/7JS9JG3glb3nmsp
QbMfkL7XChMok8tLjaRwZi1KhwHfOHxStl4Z/pvAIKJVUqZVQbE515Gogl19h+kKWZnQ5MP9ptqx
tG3zsAJjzG73yJAYeX9qMKvd2Tt5Q02XePpkEvqnBkwDLI+DK10x1GVsifN4YeI0qd78QspXkpdC
jP07sOcCQOyo4od+RiAYFoUBs8yXxG4/mMyqBBkhykIj0D3CjuL1t1s/XlN+VCoQlizar/daRs9f
205/6Q0Kmd7yzwCPRFs5Q6B539r+akWW3nXAghEzKaKTWXnw7bLzTBCVNbrG/dao/lKKG8Onrmk3
nRyhOM8QA9IY24XZHRilE+ynD/5aTi42rjL/QAHg5Cf9410KjBbpIPMIlhJr/45fm4hP2BovCITe
REA6WFkpZAD0puBsBp7yj3ICG+ybQMoe6u8KS1Sf1iDQmuGRTr06a/Fpv817z9Zjko8PhelZgFJa
DKjNnC5qu5VsoJcXuDA52zBMtCo9Rsz9PvpZdsWwATpaBY96aALDVJjMy1fTGiVZYL1rBDGwTMh/
OD62kgdjmGZMN25S4ZtTB0x8Ab/fatnunPrvPCO/HH37/Sm9knkF/7c1QnZI2hg/VLVbcwierOEW
ydQNs1V5bNvZK1HWfX7hy/IDkni8iAw+5VcwsoQigN4K9SiB8wphRdqE9qXZcOzdqyDo3J5IUh2p
NUQHfVB5/3W7h/WpuiHYpKY7W5s6if7iJApvrwWu5H9e10nrHdhZ1/S+oLx9gX8L/j114InTzvvz
EBq27Qqx6EirzoPHf+m1qKLUpWI3IhCZbDGqh80TOAr9VaJOefMxAc3nXxSQkypIi1qNXQlM7wG6
xxroVeHlqDivbSOGpgaKx97jLVIdtXQz4/zTrRPEwmeSy6mW/wzDWjqT341CHheegoez5h6mKQgJ
oTZdSxySMMfQkyRKJASfBxMmh9T8z8Kbfp4FK/auyluoLed2e40T+ODFFxO2wMApkUz3UaWR6p/X
eeBCcE6d/PlwSt7Ln91/4JPHzcNUugCeTs2oEREceA8quvzqmhx3qhURJjDVl1AxaPsH3EiFXUBy
eZPfCqV8K0Te6xbVUomzqCUoWm8dtsd3xs9DfGIhUZxl4Oy6f5X8AdB8C/T8InTaZt5+abf2ZJd1
tsyfkva4qU7VnNZxMw74DeMqs79dI3KD3rezBOtHaIn7jjGyS6Gp7yE9+FvwNMEZTvCFp1/1EMtz
qh+clq20kSMQ1H1oPfNb0aGbivaeUNrBOzgdE+aZHydp5iLAi1rFEhz4H1ZNYScrFI7HjCVlAxXW
/nfJzaZQ/EJWo5FUOjvCpPS0wPwFCMxeAlynJ1P7bLIzqrO4gWwi5nh8TaxRKqAGM3OhUDRheK0u
PmVhLWvqhfiEPLCSyEPuKHj2dpwgSj4PFMgl0wYv+akexCYkxVju75NIAlvHWnkyeX7aNNTuPJ1a
wTxgbPIg/eMgnQ1q3GDDvJksqch4E06FTRcOomOaQKsD3lPLh3V9cXS6f+cbGpyrHyWviClI8wyc
eF0gXci29C+eXx+LXDmMy/83T9dsxJozoDLFMdOq+py0WAziwtP5SkBmQMynS4hnSEI17DLmJ0Fl
mWxKhegRQUzfpQCPXt3Qqq3jkhcHV5+QWfruKjc52XToibQ7lIdAemzpnZYQZl9De+zxG/++qtz2
djeFMbWg0F1wu8zhZV+sGPpUXUe3mXvSrUMenTFyB10DRdXNyt3DfQtrIPuoiKpsMlzy30rxm/Y1
U2d6OMjIFbDDWjoPDzHVzlp74G4o+kJlimIWaEs+ZR/fduK4Njat6yWp1rPZZM8lY0BUWOCMpcfs
OdjGeFLz8JBLtoWU+46OPPsvTxIhUks8cvR7TllG5NsRYlpwJ8dqY2jXBAD83xT5GrgHnLjKVmr1
y2uwWyeXeCZaJHkCUxQavGNIiZpAJPqBMBJ9aa2Rl+0iMABiMb/omdReyHCkDYOAjnRwUaARI/TI
3SQbTDNsOosB0HaXXkp29QmWU2lPhDJzEDW9suX++UMH2HpjEKHDg5OMDwjiEWOfDf4xbzMB2/j+
GUukCA8+ermyKr3lH5Bj/AQbKgd+KlaAhkvxpaskPm6bYsR608oycM5AZXgYSg/vLpxYbywGpIhO
SqKhTvCzmygVoJNz9EHWnxNHs3oGnFMzl9H7Mr1R+0XJOm+wxUc4CJbMlROWFomuQWHg3+HnkVTE
fYJBNnNXCvUdsw0NQ6uzvesBbRJ39Hj5/pfEQPFFHekd2Ia3FqhTKM3qBjQHK/PjBmASPqFghVDk
hs1OdKfTyFAZYZ0A114VrWjJh1KPOr+Yy2cdnhtZofJ3IEIxo2YvfXXjg7OKBwsGOmLHII0kgp9d
MVXnuyC8dl3LfXWtsvGU9rBaV5SX8RfnqgjlzWUTuj1rRpM9vOE5iPAkAJrk7qwoYOil+9OVmcTy
3qAQqSPEk61AfQLa2Jg4ipk2c32XvTMOeGE2eLRGrfJUXMzCFBCLLOyMska7sc/DOmbX04ZYbalY
tNT4IdsYZwBx+YgoVsps+JLOZmzmI1uwHjUW6zM1brIM7l3ipbUk/KGWzsoK7Y6Nf5+DTqXPl2u8
OalB/VO8bRK6995lc7sibkdJimNkhW5XBbS96GMUr3ETotNKvZvx9qNbKXk/TqlDNCh6E9L/XFCU
U5D6bQqFhniWJf+WHX4E/iApzUGQdMoBcjZ9jcS/w5UbJGSYYpiR+jM0tWblVAvMX3mnIjz45/to
rpIIhAA3JYQzP4BsCFctWes7ydHCkVeJouMO0jESsMFefXxMJj7va5VSWqWI1JHCjaY5fNib6JxP
oDTC2P4/+jd3eowkgN+FXtFgP72Z6BwjtPAxLtb+b9qxPSoPhMFR921m4j8RLpx72H0kT8DAoP7J
uvmgJcY31Bvv3ibR97D7slNYteIrFaZXt1ENmk5foIRmwMerJLo2o6b0aHrRE+w46A2RvgTIhjFW
7eRlk6NqrRW8Pm25Vvdl1UkaUbMWiVm5csuJx5Daedyya+dC+/svvr2OFunmYSvJlCGpK6sIplN6
xC3uSsTFoN3ZMQ4n7rD/UBdd0G3cFQ6dKo3XMTdKaYJLt/xNqvZPv+Yj0uPlq6lhiQsyGxRECbKn
he56kJO8rApJxy49g4S7o3sWG02FunVxGs1Zg5IGbAC3TvTe93NfM/3vcEFwQbFFV/UmnQOn98Hp
QE3E5yuBq5CErYpwZVFl7NPBFC1uRS2CPb9hP8VykKq1QQlz2N2axnBylQ/m/b87yiEv2nKlu2bn
l7Yla9bQaGqfoJdiLU9qgAWvGkbWVjqV3Hcatq/CoNQLN+0GquMRipdVr9On+WtfLwWydHyRX0Vk
fxo9ezJ8ImrN9GFjfja+MjXawF0b6wiEbxzNrCWepmAQ8TyDt9PEWBFAxOUhuSd0RHg2g7ij3JXY
TISWRwP1RK5vyKA0ZTkvQ0nhUC8pxiG65Kf0Yq4RGZQ4W0y6L2rPezB1G+bhmyVRQbH9AlAYWxaj
JvJ9n9S/V8+tfO1ZeU1ii3YKlnTVmVS24/GFVOiljCC1x75RE6H8Cu+hUeDVSZkefNPMBR8xrPF4
huzpXr/EHTi80eGwbITrttfSsJUvrkRjdlp716QM3aNRMYSfpCPW1IEgwKIR0c1b603QiL+gz2pm
N1cToHpnuYI8AtT7A4I9aoaaN7puKwJB1WIhbv23wsC3OlpwTsDjc1D2UCMl1Hqze8290Uv2pK9M
VfIX8JlyahsYaZzu0bwM+wE3cGo+VVOMi5Fbx8TyR5Pty8mDP5BWojauAUlpZnHzD9vSztyBNl+j
ctnlqYwzywBKSVWKKQDsnpTGRmTaRmKqcoHyA7yLJKbi0P1DjTPi0hHJTlsHywb8QevA6Iuvobln
oGPLwpiDjiUYQDYp7wC9ih9SgKk/hZaNdFKmn9JFMc4VkWnblao0dyDwoznWaZ3ZzbcwuPcycNjJ
vuzw92EK9dHPnrlpGIZ1zI7mc9kF976u4WIQSCxpcndO8PT6tmtUCY3VyKSUoBVqoGUTctybxf6M
HAG/1GteM2yREoaQT+5iTCYRgWkIqmDi1FfxygnvXDkP6zkSZTX8jvk1Lc/7teuM0qSf5prr/2Be
CeGAROfayj2l+kCBJwaMyahkzADUKqGR1PVHo6xf64Dy8o7nBWch2Dlf0Sl1X5cHDv2E3oRh5ZXV
GcdWVT/u982JExvZZsibOpVRnqP772OvNRzNMsZZQ3WNI6Hg47c/7m/dKocmAPm/L/dELqE+FK2X
Ez6MJ4PWRMC3Blq9SsECtjDQZnoMNPkI4Ijb0zoy9dKuyj2IZOvy9UATG7Bxs05wVHYk9QTAXD+q
D2fec5Ew5QgD6MnjXJuUdZVb5aoK+WT9Yu1x4yqYKD23T3/Ulvjvv3tMaTUS7OTshamoRNz8W1AU
sjIGPU2CoynJPNJkk91fccmWm2rKIfFh2xdYQQvv3y/a6yZYDb0vwubm+8DQbjwsv0TDEWqbfVOk
BDrOb/O4gecKinCf9mMfDma2EHhBfwFonUc/gOPXMJa1OQsxOhq8eIlnoSgiwGJAB1lDV+hwmPFz
2awrbQJvEEgcXc65oGiuc9oXd6MgXtFSXWigJC5Xoe521bjgoaLgBume8HwBStpJB31Kc4g+PYyA
YDvLhDlFbWYFLWFnxU6HuEKiBymCTL81wkR13C3FFSywtuVsYB1H9rdrS7My/Wy2Xo14DXqJ26+o
mgOWlM4cup5G3RuQM9W383MBsqIS8Icn0Wqy1be9s8W7egAEsNzO96NKs+THzS+P7qfU2DYp8Y4M
Gh/kR5UPyOBbUuuZD4OB6BmyzB9MJdhQ6sF0MLZfstyAa9QPZDz2UgBga9/YYys5n4JfQJgxGLM0
A6g+wXtZS+NNpce1BQ6TjwHP+31rcOT50e/R2ZSJEVy0v2E7vFlSBz/k6e51N/Zwl9MxLzw4IQ8d
gIN+mnGxkicIzMahurb85qGMbU2uFoojZF7I6aeH4KHHK8YLhiuf5K4CIRv6TvM0khvKmujPA7UK
j+vA0ziIXGwM9g+nuUbewV8NV/KtLdLn7Fn44QzmLb7zldnqtFkgVkq6ptI7AZ5ianZexD8oDzCJ
GFfSc1nMx6jYZ4tUJAS0RO/QXoMaQNneoJwotz9xJyC1s3PHoYcsU4QwrTuxIqJAdWJTZ0fmb8lr
uJN2pybI8eh57uBLwruyUG6K4l+zxGDMF7Zy1hKLJS5bqbb5Rc8NvsYnGObNuXz11H++7gmdgjtE
mDQwoav8SC+IEigDCyET3TewXnqyJhtVoNAoNSAzOdWVWu0YyRrS6UrcV96EVr6cWNheshEl9HIq
N6TztM+tq+Hj0hnew40pYObpa6IoGZ9kvpknS8V7VcySI7ZOelVw6eDh7ZeTbDLItv9mElez4Lj8
6RM8RsWs83S855bXJR6lVvJ41RZiruf8+7zVy9A5i5KsEf5IXlI/OitCz4XZ4e5BYNxifvRFoX3F
xbi3o1cU/X9xC8qMFAwcVCY5Qt0E98de5cNp/06UfpmJB5DdKmRFhSJaPtcyCumjDo1vk/krQ6n/
myG5PF+qoVBexbGdc0HCTFfjWpqQOaXBSy3u2ykaxVUYg3Kx/VZ+E83ecAiJdyQ4/MQIWs7zbhWj
B9L4c3ThvG3uiNbW++BDHUv4+zYflt0tBEiGmlVXpsBXvXgLjsxM8QY7L/NtxTZFc5zcXkcYeEwt
S2kUD+2mHhxyWwAzFXoM+Gqfw3ooIsm7KF0D9+fduI37OJOkmTIDNjIO3TULhxi813nKVGDBxt5a
fQWqZfztLgPafjxOMJpRy5nrWrKJ14/rk96P/knSVNbqfmoiZmRyzbUg+kh194J0SPwJ3pD+K6Js
MHpHW70CtEyLVVVBhYfkEcZUqGIeTGZQ2/yUlSYF21YVsoRSrqnCZiWkccpBa8QboKypSUiF2zeQ
P4ODeuH0ip+UpBaVxDnIkIf9/g0zpJ01PvbcaDG4AwK894p6G92+o9lt0cZLiJo0LmvYKo3n5ijP
2rzJqKZbe+6RVhFvMOQ9noWlqNujBwo2vrdpWilL/EE/nduUhM4vc2cuE8qZhXzYD8u7RA7DLubG
3geKO65yPyvvz+s6TG1pUodB7BYH+Z6BngpAMDipPBh3545EKvcBlTPcXMkzqrOyMHFMDNcKHczl
Cj3p7tj61sSYuY3lfWRmo4zkHRTYwk8Ay2y8y0hTc69//b330weyH3b/9ezRuR2ZnKEDDupYdlnx
MxI7JD5CvzlICxSKAURaENP8918utg3hWRZd07ipHe1I2I/SpqoFvAz+XrdBhj+esJHYLGkVrDoT
3Cq2nw8yhIholOcdBBeMgYjdydpFDhlPkcUhx/7NZ9sCTUCEDRXc/LTYUlufph5gE3zpDTpBRGb6
aQw6Y4Ypo/jNpwjp6AiurVW5tYGVeUqBjUiBGdCj6Ipoi3m2pvhczOp1CAvwufqLPXXRMlYmaM9B
bPrXpQqXPkzDozcimaihw95buIKuK1clL9weC/WVYO5UdXEsOYcBk1PlNh0zPZg73mO9dvyZnfa8
tw7BraELxNQOA366p4Mm6mUknbgAZ080LUE2kzn0o4wRjhO4prRlF0vq2WXUpDSO6CDssc3DX96d
xVEY1HNt5HeIv9QhT2vWdokCkl1jB9YKH8jFhHrrY1V4RznpCzNvWCdTmqc0YiBFWQHCXFKiTA+Z
zYVcmWP6LpOLs4BCVyaoHOP1H5jKrHdRhh+2ZDth5/2pzQTdOiKWF8Aq3XuEOgeGpsAgnSyR+29h
N9ZP0KcBZK6LT4qQP9b6iF2/xuqoOqvR6bXaGDcG7b3UxvlvpUdLyyk7yVd0sD7wgYTQaDuJYsSL
didXHerQ5qOLZ50fWSY+jndX4UaoRKDKCjW/bYcxGZTkMhwEDVoCZLAHbJPI7nFkxCfsEr0wfj2C
XVmx6q6FsEk4/fUyV/oseHHX2VqOY0qPNP1Y4a7oEJWjRZ98z7IxPN4XRJQa1JpBuZ9D2su5Kt+l
KogUKd9IGSHP+K5120C1ASukIfeiBNHdyUs6k0fYEqMGAKDVHVOzI9O5Oq0kaRfYMoN69mwQk1nu
zjQhgH6t65QibcYUVIp+0t0I0e4flPL1s2RF4+FxiUAwUexJSkA1lts7i2mPVmRmxV6z5XEgDgWL
0xQDYptIWsjq/UBo9E9V+4UchTSim3vrceoVgTcEScQMXabfUtnwyQJazKDRIZWj3IpRjFJ9oAOp
fnWMTgHmfWuUcTBwT/WfEsJBlTkbQypiuS8v/15XIi2jpA+TZTAxDuwi4Hurs9PvZtOOFU3apnUf
y4pchfBIlK+YcojDNQ/mi22LI3ynJzeuid7fjMST4TZizeKwJizXHX+dsA0VpllOx4fNfJk6mXnA
/aTtV3nt1paao7xP0VZia6EGnAYSi1M8Q7PcV4q0A/ctoQaC1aIxM6fHuIuDDIVlJIYoHQt7ljtm
+EMlWK93DL79X6aR++DjV4ez7pcglC0yrEjyWoj9HvNOTURqkTyJ1+7rpemZe28xuojxC3eRwhpI
8NUlsR94Vx3OzeVM4dAPjuTpzRIhJiKuu0/4RDA9Ju8Fxe/BevOnoMPE1h5qlq6wcdQWrgYRG+Z0
yBtpkOvoPuZ7hCqi5Fp9y5cIrB9SdE1yANIHorbsyMzIW6tugCd9pM5UycjPuP2J3Wl0XTD7qS+Z
RrNXSZUfnWMNtcxvlu0vd9rp1Uv7MyoE/slJVBuyRMze/tMwXSm0GamDOzU5pECUeGsZ4pRNicmc
wgoXtjUljR27xRHthQTHS9R1W/DV0O5Wpz2IduqynUF7LLUHaruH3QUPMGCbwaRM4e56aiDPpQTw
pyYxpxtDWxmiaoF0CJ1LuR52Ry2yNhD/Q2SbX/XC5S2bpJoBEClQzAnlcc1EaHYZ3W0XgGeC6PVr
ZruFndSoh4gCgIGjjbBgVLlUYHL/dVflviYGtpvJErQMBUsvJC3kPfIYKEtsZvS2oweJlgxxRUQU
40z+5IaHA1oFBB7XfwG/PgSIerqA2XQgYejnjmQ4azP3w7lfcMJ/nV/FBElg0i9feKt5QoZUXhgp
OG5GR1vlkwpSxEX0X1yi3X/nKCiSem0VXqjiMEAb6yyTW95gIHr9YuokulqAWP7hdQPWK4sv6/VK
iH2TP/00rMcdljF0fx0tCu32PQ34tw8BxODPnCfe6h48iiHHMEXMww2h/fKuGIbnze4n5KNaZu4L
nb5/VeDBQ6zkLTiTW2ouzL9IpIrraMtoGrJo5LKH9bY2PhsmJf9uF3R6wjYMdmwKPCxgqFFGtQvz
IsUsWENQOeq3u/WOdH6dLNmUeC7F4Rv0X0svZJMFFNIDPr2GaWdlA857XCbEVPEgi9pfN7UzHoy3
ofpY4qEs7Jq5f9CxVIkQYffzi6oAOzbYjPtjCWl3FteXexIdm3mzmixNEgnVY63BPf2pWg02hA/+
WT/IkTFr88PFBEp6GeG4UKAQyyH+ve1hKwa0xtMlCzYu10pvh8RLKXgEpCbujxbEH8x4KAZsW0C/
NKz6FYuPQLxxaVpoJ6OQhVkzkTlOEEFen/TJuSKaZKp+D8xopdYO6hL3GCHH3nYP9k0CVy7tAqC/
KOa2ap1Ruoomp+bHoXfP/Eb4tC0YgI6XyaPiZByHL4S6aU49nRnO1b+rM3nUJXgyIizfShls7T7h
cdn3krANsgAl/ubPRhTOgbjYRcg6/HaH1QjxSEM/loR6N8R8f2xuikDXPtidCTJ99RxxB3EIgYvb
ZLnSXTouHlcMhDyZnGocc0ip1RvuOjXTYotpZLFqBHffifnZC4N/iRceC58yXSkwk8xdd48juQ1C
8rJXi9xQ8SdRqaRiOHpdMeUUCWAp4h8AR2bzU3biyAiZ97Ifi8oAt41xQOBCIkMuGsCT4JwyXayw
6756ppBPYHxclI9qyYUPXHUw5aZHM4IjNm0TTyjnGaWApz7IOB2G/S1Fpf0/+1uV51AJnIRlOH58
ozc+uuTw4Lh/KNBvxKBkMggFmWMmD0g9+1FmA2DX5S9O06dg7Agm921hatEF8xjK83XcgdK+fQq/
oSgS49Qe4bh+it9hwTNv7HJmFgRvGfQxRArpEiKwzSTNOVHDf5dEPILK1fLuGk/4Pp7S1UoiYjkF
Hfj4yk2FE101dUjPrZItAS5F2z/8oQc4S6MTV6kfbLHxMFm09uNxyZTjR0ofwXwgpbcH3capM6pE
lQTU8nnpqBTVQ+Zon6GApMzLNif+tnuZSPOJy2S9YpNrZe8qLXleMyAWxeAMmWs9VGYnmWdv/v/Y
JklG0AAsYXUyqM2w45mfUZp3fxE1t2lJlZzzkUzst+8YUQwiR3LY5gtG55Yip2ahfB60kW2Lk6zd
0U6Wco4KvkRLpbwZGHKKWa9+CiWT/6fO/Lk3Rjvs69AO7IZLamUFMF/UVDSkit/hbH5MxqoVewvh
i0ixjngPqsPrCsd/6wJJcNcRrdsSBGhlnminp5zdc/kbGnitQCw/WEoFM9OTrv6LZHXYWGh/z3P7
PjLtaO7LkhPQk1BhKyV7533ii6scG2H7CatP+R0jpo0iP0Z675qaBw/xlVyzse+SHElqId5flIH5
1bS2ajPkfBP6sikDy3rCNQ7i5GLyASDLh9LvXLzvVQtYr41DwAKSqWoMzXGba6ovVGJJOpEOF3NJ
VOO6+xSRT7oqMj140V+L1I5dQIRz2rzQqXQlWO01sNO0WevC6Q2SV1rHZpxs1nAZA3Q46USxE+w0
4zOAyCwHJWxKU3deNJ9Tbru2m/sxeTb3+Kf2ozi32Pb1y/zddR83o3TrZVgTkkZe0AREwGm4ZQOy
jn+pl7LIAMBi+GqgThEAg9OsrO86po9C6vaotMeg1dyegtXDxxMN7804jfKStNNhXAbn/XOBxjm/
M0YoWMxbeGpWPyu6kGrKkAolWI7bEAEEEzuFK6H5GbCLCrhuPknVvKQpDDYbFYp3ua3oIq1UTnds
D1hS14Ch4tvm2zGVrH2oiARjlZKGi1dAWsI8z2YPqF3NrFRtIO2dKs3UEIlsnUhYCZ+PtPdIzXVx
VhnzIOFQZN5j3BlKVhTxZ27F4BS25oHQsvyO9DvMom1rLCOo+sSOn6VA2icK+RyyjTmPu5jjo2q/
aI1sNw3vOZFcy2AGBD/vk6ugQeuAAYy8/MAZdGiFnW+bwKL61RHS558FJ8EYAhgO6imwgLYtnxk+
xilMoXO+HOKCYAJakxB8UObqqbHMSwXHvf6QTqeE1sT5gdvTBGhUSPSjWzv/ycaczcQ7Wmrhaao6
+ya8M76eXgljOFcsRn6m/x4bfCBoMoILZvrqAgY2oxM+BI2ecc2WW1xcjbjI+z424WX2kJW2e+BO
DpL9AQo5498Lj10EjOukA0aT6nN+C59R338a8BWdcbxkUzE9rCJopdnXCaMnxsky27AhcjMcLq/1
LlPtVQDzJY/TEsIOWcty4E3krMA39bMAcaC2BGLIvtGc8PJ/qOMKshwZ1S5MtOdfjDogIpZjgyCj
SUcbR2rbwiEEojfHhe22eSwiNlxO6aLkewSUrZackgrGh+GRdRIfje3qFkPtXRxvqP/p7A+WWWY4
diGnapZKvJ1Je6Ipp+JxLqAbfDNIVyrGMJ9lS/7VbgmJn33UwBQ7sSrHRE4TP60G5YsLhO6haPeB
RMuZdAS2DWzY55HaGWsBQM1a9bxlCU1tKMxSXiHMJzm6N29DxontA90vFNW2PE5PpfVkSfZBBayJ
3LaYh9sicvsKP7752ZDiBVpIrmO95VXf3PpP7QWSSMIPVWuL+IH4tsFN0SwEpeAivQIR3saxA5vE
v24eilIU1fRKOY2KqRWC/iN0PIzbE3UM0Lvmk+6s4SgSKHHc1o6Me1XeRRFnWsIx9BroBqm3VX1y
Nh9uPXst6vLVMh13nQpckKufNbqtQ0u2xSrxFr8trXGOFUmnY8V1bAcOpsVU2np0H2fWgMoHf+XG
gGLvv8we2j3Ng0ijYYoQlDizphDd5V1PpeHje0jbr0O3OvefOTUNlh254bfT5VWWKadyUp5/N60i
mkEB/3qDSPnLMoJziP2byoP5wWNYWAZf+hydssvx3Fg8Fn/8cqA4iKMb45VJu5BVxdKepALG/mxm
Q78v80D2KsYJSQst5p2u6dn7e8SBtShbSc89kFzo4WoowqUaWICkET9F1Fe5wkTwtUrQSHnlfUHm
yC0sY0jqdK6nCI4P0VI0gYhhaQ3bWIOBoAtZnztk3exqj0wA6NtEFE8I/SZ6Y8RfwpfYEuNx+tRJ
+nVsngfDE30hkBEcEHGavQ6aQ/Na44cXMVjpjGqOI/EocCUIWO+nNQFrd+qTQsdrWDn9nhoRErcf
RjcuUpx31xlvIaQjzXIWNZVukiqzw6rKWHxghAFcZv7ZSYmX5N7rSeu2V0mmJg4idCL0uFFwfTGD
gukakvA5/cupqlWxtmUZzSvyeDfhnImf/QutHHTmBUM6VsbUC/wmINYn7bY6sMAvnlGJlamTdBJh
e1NndAeoGI7Meeij4baQeBkfVxWs0qaW9TGRaFsK/HL03s9QR0E1gLbL/dU2+R4ZOtirYwKIfiEX
dXipBwefP1KvsN24L9TxNRM1qlEtVGBFGMl0dSplWuBxukl0lP01vl0VE1crt2pO6SviX1wJc9kp
uwOmsm4jrmXK8bsphzMP7BcJBu/4t+so2Rw6XBLfExonDscNfc0eAgurIIcX63JtVAiBPtWr27/P
5HsOwKA6KhcDzDg/aQIC9ZIZ5jJ9R6xww5v1IvqF1DnuAwMwdvQedH94pzLKyQ0oog95yuz4yZgM
5EVEDp5QYgFlfsD1xsH1L2ONf6LuARYV+NRGvXdGqsemiJlod52w86/uY5ZbI/byJAsWtgg+3Jkf
M5vUioxhFGVcZ20k51HoYDZgk+Ecp8P9JIoNUcaXpmPNNfvFCli9iWnjcftrQkHSEyfglD+kmmp+
fosgSk7mrFgZpT8lFi+f/JyjulWNWnxI/iZZAh2coYvIyTMT9oSg7eB/mjVCL950Rdg8YjH4fQnn
pJSzsk5gc2ILz+y8mGi8GHJLqeg3d50del8NzUXYJ36Ql3fud71FWaDsZw5Uq+gclsrBA8wSucUO
g5aP9WqFCb+gnY1xYmeCN5lkKv61TOZhRmKkjBOR2KXW9jla8QD6cNuKRQSavab/w+JDg/XspLEO
nXhRkww1P5WKj+DE/VMNgl3Q+bpjg2yN+d1GFSrPCZcn7R7Z/Duuo2vszEYnKzyYCz5ATk0izS+E
85UqOZyteeU/9ve87F71RYT4i9knnPUF5OhaHSUsKgunSwyymZyR7asJ7yboIneMBLQ2sVN5F+Qb
ELoovX94WQwYbX4OU3UJsuB7vLCseyQQIzf7Nk6/sL8KsJUZkOPj9txVNLqf3rh/ghjdbMpdlyVW
UnG8lLPwQvFP6ihGD4OIaPaGagcBlwQMFbAWsLdvnkODK4MTFfPwfj4754WbByQnElGJktsVYv2H
ro129fyUsKfUhi7ycasPLpz1eXh+HwmK1CadQd19jUxxgk3j6LHwYmr09Cq6thPrggei7ZTmrl/q
ZAPXHr7yClAs7llX7iNFTKsQwbEfuh982k4p3xgTncYvmHCqu+Cabn2yCUUTAGs1gZnLh6/8kDhW
y2tvD2/VH13klSOqHvWsQof9RoS+JFCVV2cLghgBaT80B9GHHL+wLPE3zRiYuYcuDGfpXc8us8Rd
NeaSjsAuoqsJwTBab8UQT44V9Mr+U7NYl1+i50OgPMSIrSf3EXKsZ4JwBwpP9KwYcN96YI3sJJUD
cEZUgLiZRJ+KzoYFnJnF0bYXMD5vpb/Bm5UFBdeKcXJrfqKWLFqIZxeJ/4ff81/0k1VHM4MlagsF
9QuKIchCj6zCkEYbhw43xiH90xU17goqwpUi8i2lM4qefUA9qm5IHN6uRFwQQT5WkXd7HDFVCDoq
a/9R33BBm9JFlhUp35T35avuLz3SlT8zyl0ixmHIab2AZdhdK5h8t12QlLY38bNFw/55y2VJbXQQ
4tzNwVvWd//fgcC7tOi5KASVPHmfg5Wmwk333kLYjZD66B3FKuIsk2Xy52JxiipG2PEj5msvUo+B
xteSduriavY1EqekbjUv3aix7fAdk1qWfYHtKKHQ4waA179FqpqtKsRIhn/nMZDDbLXVB1FowlCz
I37hmPHpDxpS+H2eCZwfxZBJqLxHeykmcAhGCMkOpbXIbwlt6NmxCddcRJAF3h7q+Ah6RS2M1zat
08hEHbzRetXUQcevTKo6U+tJd35otBWQ5Puugqz+OUPNYmnoRaZ7oI0xYnqJcQRZYGD3LNSAOJLt
WCsQrvIG7YiaNCyIb9TMFpwISW7f7SaoAMPoUXqv2wOfRrKG6PbyzYY3Lyo2qu1A8iH48E8sMmsT
QhEb2Zw796j4FPQgMdDvWQiIS6jD8UAB5MpiTWxciQCD/ZtCT38uWBEHsXmikKUh6Vc+//DLDam/
2E2KGYIL0zvzo32J9hShOiaU6F3RFb3UMQKTRWx/L1jFJsqAdMYwpR0az7I2bLmjGs1/g3MswMvn
zDXxkeH+MxrjY/047N30lnarpumvCDntMQQP3xz03U1rj9oM78fpLfuj99XD9/getjvunBDcDE2d
cr0JHfF1Saq9LTdPHvcpEM+SwFmcv/hqnC/7Kux+3oo+L1T4oYKcu40qUP8Oom897NIroJKY2Wsz
vuG9UJoHJjejO+YyQ7T6TCIfHbcISwqIVBVa7FIrPvj9w1wS3yW3Bri+kDxCxZ50G6UKIZYcBqSf
rAMuni5BwXoSeEypUOhjlazooa2Q3nIjhuFhVMjBdysBiUFhxDqSdRK7gSbr56VBO0oCESfUC/O6
ZmY6UdsHI/mbppt7EL0qUier8bZzkxhZn3uOjEn2bg+TW6pUGqOKoXWZ82Q+pPuJAI9vIA7TTpUa
+4MW2ab1LAhsqjhhlbeqbZTzX6U5v8ji+lbZsThdLc+DR5XszriHeT+uh+cuti6C+rU7r7yvKwwu
bmipMx8DTniz1uhlHNYO8iNHex6D/Zsu5g34GLlk2iuFEbCszjqj+x8XvRC0DUKb/ra92Y1Kx8Pb
nobBnta771SRzCShWWxwdH2ISSuLqn/x4l+x+WOp/TAfOmWlQhhc1/QdDunkU1uypBwYdQj4NzTa
d/XC2hSpUfJmlfV4L3DobRAB+/oiWQhCYd+w2z53kNbt09rps/QQSx2+oeczCnc9xPD4LjUm4zTF
9OnaO8GKHsL0Lw7NfRm3VkJEubeUtgrfsr5TxBOs42KY7OquAUD/E0irZU3OEXp5v6xMrgRYNLYV
YK8rKJHr8cyz1yeP9AZU3IEOEUJtagTqaze8ChVW9EQOdBJWckIx5RDuLmTJRZTf9hrc8nwXEmun
ef3hul3jckmZuLchV1RF6l2ovhdzus0dKl9e6iM2lfxlDfjJoLgpAPZk0ezBRs2idBRQ0fDqcJsP
UVrBIR/R+rgSZWAcl9HgVB4hlyv2b9G1UNpQA7onBNHLed5+OY18Y7OUtN11rLdqrH27bKXcNKVT
23Ocr2812kR8/76R6Q4UQAf8ascOaThYUlqUmfyHpz9kO2lT6Hi2ixdp0XHrZDOFxawNRszIAnuS
ze1nqbvjuhaSxFUmQRlG3jH0S6Z7ZQX9wTDW0rV0q7On6jM6mSjAwiEApauMGbEV908BzYrxiyGf
UaYHjPjgyUmu83/CRR1gO9D9CAxeq5z6UER0hVWp3bP+X3oc11Kvg+vYjUevR6yfVh4PFXLAFrlW
QK2N++ZY7VDgPRCRZ/vYcG1ssRXO3DFFqdmj0z8/Rq4ixTINjlMHw0hqfs86UTIArf/5hFWHtTAh
qC5ZDAKWAGqQwLd2awgCzdSk+Gde7bGjRIAO5JjNKBzL5ChelGMQzV+3u03PSWGtkgHalLuTa2sW
FfeeTNAxrIKrHaawvh7eMnbGU8RI2673Cf3zwA78ROnImbUHO5CD+y6Z9TVL2+Ae4/iGI4qfEOZP
nadCJmva/gXkbfRpB5UMtKIB/VAC+20wSwmI+e0fkj062dxUp25ib00pmUoDEyTOikAsLCbEzWgh
HP0hT7sWvuxFIZzjQVl+Shwj5pc2MPf2e9cdG7dzOtjt1rf1w7QGQS/Sf82Sh3kLxTySpha88vJr
afp0vryelKP1O/zmwSq04GStWSjwq1GTySRXSHrrSF9Boqx3p51M+6Z3v1mA6yIN/FNSNyOzqCL6
XmXiWIr0vSAjeBNIufApx/u24L9jJANHB9eSIUudnjnw2JkcAif/2yC56kaP37QCchATTt/U6ygi
ArzkF24nHn3uAGgmRFef5bu8mjzQvVeW47SFwf3DYhGUva7mRG+jcVjGTMAXvfvTUmzVsp/LkoJP
6H8PtlEiab8t+br0xh1UXes7WoGkXokpZ2FfCHgfdxTLD4ZyXBFwtdZa0vwGg+aXwl08FzIv++Vu
gwy62UPQsmKJuuVmL7ObNqdlaLkgmOGZez03B8EC1r1o3/kM3NjB1U+liU/ze7pFTkL9HVDTprn+
UFrvkY7SrFXeJWFjbPGKd3F8eSTb5rvkWWsfjb8lPqxOce4mNuJGJQOsp6wcoX1zCc/YWcUJZ+b0
4XfTgnJWN8FLPVjkjAH7kYesWKutk9gdf7IG+g4A669hSsj8KQVpFxuklIoqpgu+TBIauoSpB42c
mn4gfoMCEMtAwQA9oVp3EzqaLfkDFAcd013LI3LKyA15ry6j3KvvhiuEz72tuewIZ71j2lqxhEW9
li14rDZK8m/QWJnQ2uLhbH4WPQ7h6/IP+CWFbEmDjOlj+f4RBlanOaQCgwIwoDekTb6g7fevnZc0
uTmi5PSi5tEK7Gh+TeIzD985jxzdohA9/Zo0LuO+uSEZTNkgqd3MCHEwNgInHZe+aYMgVzFthXmx
edTuel5HIZ+jGzt8RsEbglpgyYXZ+C6y6NSBFFIK3W41InUbYvdsHapslcT4xcCRs9CzmMhctt2s
jFuKh/6h4DZtq9XP0xuh4uBCIcrnul/52SdfOG7x9PdTE8fXVcutsXlUbNrI/VjA45nQPVa53tQ0
NyJ8EKTLcWwd/ldUEiRn2LzgC+v9Ok/YUKmqNzjXHOqJIFsMil+cNNQw4u+gv67mV4vxGLn6f9Zi
wr9WRJnFSOrw/9769XLHWBCBwaJ4A91reprpZM+a+s1/IFMIhX4YH5AaQ70vecu4yfo3icmD5HuN
RXBGMsijNGRQD3x7YQx80PzF1LnSqNP9Tg2WKurprXSq5MSVJ9F+TMQZWaC4MP9TW0pY3uh8sYjG
BkjTaFfBOe+Vigvo0q+apOn/JIw5jcekrfAXkp4atcIYofq5RKotatZOXJUnMXH9VEWcQbyyPU8q
f3wUDeHVCmE1eC6GVdqU8PxfW8oi7fNyXbZeyPtS9qd1ETRpG+O0yfRaN/Yvg0kw4We0OA+sW8Np
IBN3MjLgzg7ZTpUtCuNe1sQ9owmGvk/EcTZ7ORJMjsimdbrEns3iqBN9nYhGRiGvTHCo8vigvuGg
C6zrFaOtltoTgvSFlFdIzit38+yqJZqfKDsXbNUtHBhoAcgTI+PRSKzUGJGXV+fX3WCGSTwp/KCq
5yphELR/39PhvB+xeF2eblPDCJsjcx8tSHFCSfcYBw41YbC2Ricf/xkkx2en+/7s1OXckSGgKjyW
daQqsulA1av815TVrX7GJ/hsJ5llHlIzCqAnybb8LJbUSLtr5umrRb6IghZK4ThV5jxSuh4QaCoc
+NDeWAaKjYMHFOWopDV9N7MlfKspgooTf6W2EW1hLUqw38tR7UTweoeYJlMtyP+rbm1zZ9P7faxp
Ehm8AkDYu0y0BT21o5s7irtqMuG7r4xIpXcpkdxhhifsb9NyHKiY20ismoOTdUV5ZghvbEvGrgGv
zMPWqAaESYBWU4AUzLTmDAKO4/bOfaggmR5U2523XuctzaNCMzscAfuacoA/to6S2dSC9fEualLw
1LatBFfmWkwub1psZC/UbZLQUFPSwIbafXB2tqaSpjMoG/e/zFrq/MpH+0NPNhn2ZSiOuk2i1NUp
rs2qthA35Mbt79rzpbnjkuy6rfoYMx/q8UnLLfrG67yZmfcdIGPrrr21qEwHuKV5oKGArXOmoVBl
sAbybXzcz09HooowX/4yFQobM44Xjn8mRHOE+GDMaCiiLy02OYQ8K+J0v8S8PLugqnI968lno8PI
iK9sV5XKk+uFfTJ2oyt7+ZcASnOqCmyrWa1RRERDgeJD/nY99N0SwKeijGwMEdgba7icygnJ7m+e
eV2k2AjM6rMuyiR+NfGr+u/3YkZ8MvDjl3E8mq34EMAidruqFn61ZJWwyNR52TsTaKFexF3XVMlS
GZ1CB5SBVe8n7WY2CnwcVnBVkdsyOTCH/jzDPfXwKSOaNlgP2D1HPiNnlM0u1Ygyfo7MSHiB4fAW
g6hyubxygMoni0mvXifx69rXYlfs3OcJUl5Fxm3ZWVNWPCBMsrJUNh88cvwrlJM3evH9XXGfeuC4
am/pIbsVCU8RN8zH1pO0V/TRuphzAOnbgzvYyP0sCb3U8uLPwPHQRyqPmdBrjD68k3Ctz3hKJkSK
X+tMEe7s6ash4hnKCrKhcJm0vjUWqK5lhv/IyiC2fqlZSXkhCqSFgfRSWSC+HSqEhwDMYtJY1Z69
o0LbVcm0zjDmPLUL2xbayTZ3eklrmcKAS8TrnUpAnnSer5qfoz5Wq49qgQt9C0z47H3mDf41e3Pl
o+aneea73bpMpcV43tzd4dtRH1NGliJXzMm3k0D+8w3pzHt3080wuVMlMTW/I9xR1LztZ9DGG4t0
rFBqSEVPr/G2/fPLHE/1nyaWiz5PEKqpcHkragXfQI16d3gDZvhYy8417Gp+gu1QMkIubw/uDbJu
7T/hESPACnM8cydB1Eiw8g7RdN8Gnv5q9OjF1v2jiTmBd6KyryHKJTPAFZmEuwUGBDJ3DAAReGHy
mrq/0lyq8GN0LOfcABHi7UWi24HRaFRgEaLxv6BoVURi+wWzCBzw+a+Uz/eWxofXU2Q5EX1uSWYi
DrAxAnpkDaeItXuxrnHFlbPkE0nJFX8iMV6g5YBKla6znu57praCFZVyzqtYkJjgaNmC9sZR50nI
4Rja2nyWGt38qZJH7fwNo6o1aiDhbCJ9qI+2ppEeLJ+eEZ7wHIWiEwai+Nztsgmi5k1KTgrqwHPp
y/p1FmXVNJMQfvN/jgBDfLT0EnHziM/vr4UvOOMddL1SGC4kTxRrmcFKkMB7EHvqT5ubT47e72Rz
J6EchWYQNy6oUZA8ZwA2vmURMI2QDgM5io8dQR6qlLSGe5mRd/HOJtbLy4xZOsLsHPji4rTJzPTc
Ex22iAww9X1ySxNyraxRMSGrvV4sgEeXcLWJBccVxdVREAQSjFrAOaUNQ3O1WFVdkcBZ9OIwWRRe
nzdJsLR+F+yhWbUL/jIhUl65XAuV7Rj/HoZvB0EQtNyfRYd3HM+Ruo8E0sZ90S6NgSDxrv7B3OI7
5St64KIIVQ9PT4pzaV1pbus/m57foU6YHjsjGm/9pmpdnKnjO/9iZOoy3l0SGgNjS5HOc+RM/zQO
CUIKrQ3FdA1LCFL0lJZRHBQoNs3sMsH06SfSW6mJAxRSPy1o9BcbxZJOYv9vkUl+LU7FmtvfmqVf
W2pDo6lBhsjlFoSqTc9lKH+060DnBC9oWUkK/Kv7otptZfYVTKrjdRDwvkOLo9b3DOpvMMVmjLsn
Ykd4EZzWkalLnw1Y0el9PbB6tReq9Arbl5CzVtkeHjeIY1Ale712OoaTkhRo4vUL7sq+TjUvaReE
xrD4/D3c9pXowhexEg3MOsyS7piMdzZT+wJBsH9u4vKsN6B+TNsHBENfUI16OC4ZD5VJhP/0t/nn
DUcb5jQHMCvVD4zTPrniioP/JpZmXwZZbdagR8DSRRo/bJ2ofB/Hs1Gyq1xFTbBMwLb2jtZ9HKiU
BvGj3FaGI4ajHjzuD/HBMM6o5Fmd2AlIIcJ2iQ2zXQNhGl8Xs1qsbbko+sjxqx3ogF0V8mjLecF+
bCXa6TRaeKyWXPoNolVmcDLjewW5HPijW00uECVwmLDnQW5zJncb7psWrunyQe7J+7mMeBom46/Y
ZnLOyYec6l7tuxKeGjeWOfviMJX1Akx1GhQC/FF6/kYV4Alr4/qiIILgjsoP5O7SvfjAbgYKI0fk
ozl0pBwRuz+FXaAZJWsAeUdHsyktuK3qBWAQKG5KKR2RWuRbmJH2mgJPFMzJN+3Vg9cCLnfZiCf9
Mp/tcBf35xQDY/bqhHwaA6+yHwzbTAEgf4PCvZaGtr1weZMN5W9NgoD429Z3oFfxJQaSFnAPD7u/
BQKHXEjEVSdTdVdR5WVGZ5RiecpJEwjsv2ygnbdiimUXYaKrTc33LaZTSYFiLlri6pRw7G7I3zBP
GOK4d+KRVQqM3hJwpVKKgt952efHfL9WteDoJfreBtoKYoD/iZHPrt94UWsytNdQLPB6AGWqnc4W
uET1J4nlD4IeJtW4JUKq9wBx4Z0Cf5MijM3fJbhAij9xmxMuCGBGUpdsMG9AJRreSyXK/doexis2
FvWmb0pA3shkoQRa9MdGAqtI56w+OhOOUX1rflHFara0VxNtkQAW7eMhQfQm1VUoiu1v3I4gynGG
pRtQYRulYy87y276X8omSLvynX1Aa40JRbVtnzIZCTWb4v2UYBi2CYLuZPjler1SQSYuBNkPSTm+
rFgcZZzzfLS3mKfqipETPdZPHb9RNz3BOYY6DfH07ZUAumUBGX81arW3d9+8QJUgAv/kNnIfoGS2
MLmZAiQTO3mwsmMTnRo862h2/r25LjXNvKj9G/XMSZwa8X1hGmZIdDAcW2FP3fsZ75DoZNzcF1T8
aEmOg6IzCYaHNI+2xNh6mE27idbWYoPnF1xLu8htNelwd+QY4x60aoOlio9zTc8F/wvN7ML5QTCM
SIKnQMS4X5uKPuGihkbL2sVn1QbjqhelzkmQm9qEjenxexg53CeDVYQYTHr/2qEPlwLIe+Hf7Rek
r8fACOjlJ1fG8u+JH0/+Nz47B6YXk+/EjQTUku+H3IRVQtCuC/QS4YXnPE5m+OxH6+o+dFVOft3L
zcEz2qt5IVlEIg7mJAKSBbnKZUu0SNyt29zIBUSIutYgVWzE2E7FVVFDS2LtgzWvU5bmo7V7Tu1o
c1lS+ATQedEtKYW4WEkF8oiXYV6VHw96QRumUkGhFImX77u3voc9tCl1de1H3a2FdLYCGHkXS6ZS
Qm6SThUnItxoah7EydEoExwQsrLKozUKfo9oqH9l7MWqM4Nc5KcIVOx6mCnAFSvFLiGz76i0MQEy
orsfVbTIiHFOnz7nXLJK2cw8/We5TRZfkUIIFoodOy361F28t0QZ92d3FZrtoU34ADfKF+NQIbbG
yibPUpmJCVTVcwZZ30nKuyeaG1WnytuDOw4wdEanqbGdrXAQ3jEk6Cfi50pDUywzNhBV+umRO53G
CvPsMFofbsgFgIUKr26HXfKrT/pje/h5kfCj35zADSQlA0eifWMsPRFKobgpNEcVv1UzYVoBQU/G
/CnOxqKiw85qcD6AgeUX1/eyAVNKcK4Rvs+KDKU78Ju4RDphS3fs/yamSWdtHgeOrrO4/Jxq6hvK
ign1RdghymqMn9o/+SzYiGHeyb7g0vdMF+gJc0KN7pTOSHALKAWVJ8LaRhf3Txi9pewsfaVEqNGh
/e9euxUL6UM/MYQqOWZNnHBbRJqFsNTkxTtmcOOwrMCAQEgdYSd49uoYGVkWK/CGeklciJWUi58J
hYdNKROkXJzw1I1BPsCZ5Wx4XsgbtVneC8dhpdgpzl8fMzM5EB9PdaeGPuiMxWAI5/98oD0VD7ac
xx4y0wVXaG2gflncRoIrQj7Hr4n9L3Z+A3MyUyJF8EDZFSpaAaPZlkgMSkLRgoyK1Bf8EIGiumH6
WiwyDvxaxSIuOuVyTf5AvSSn/WbaG7lG7J4IbUo1ihFIsF83M+7o3wuyd9Osh9YxXegH3J5iNBoD
UKnD0BqsMRPvf/vrgD5GFzyAiQs6TVES1EFu8yIOx4tlbp7E9ciZpNUUj6ZzBUsDrLFyZrNKVlwh
qCiSy0yHF4O2R4Jv6t96dI+Ndh0GHmJvUTbWIoqWu8KFqzu5Bpp6GrQuMZuo4PATWcsoN/nLUbNY
kBNus5RdIoWnHLyfzOgiVRZR+Ik5KYXQXnnwV9rIikgospw/V30G0MuiacAY4UrBQw4TWZGEy0os
KW0DkUSJ6Ygln4jI6W520HqMuMYYaeFdVjwhL2VkCU7pI1ovQJnkcYXwjjY1y2FKQiqZncK5cQWH
7ZUL5ugBgvZlqW2zKFH0iYnLjgrVKZ0aQeE1aKWEW4BpZ5/dtcCimQu5pE9Wl4xrqBnp3xHGdoZC
u+7SaaRkpJrmnDjD3EIueMpJ6kXoYas3xTU/vS48fHZ+DaqgKE8A/N88ErDvuoeXtRxi15afOV5w
WNmFF4ZDhPv6Z8ijwEgSHSINYLeDPONddsKpXs7JxlZhC87zo7dSc62vqe/LvZ4vipFCxPvoUqVo
cYAukamCPYloleYK0HuiBmYnxNf2ZEXomSQYJ+6fm4ntjg0aHqMEbTe8IPTfEPJ2ZuSUupi8d/8J
JSEIRJUyqWWdp5Ao9ZhW9rKI2qGYcwt/unhb9Az7nREIMuxFL/gw3U03NLioFGW9EfDtLi7c0XvY
qjzYRWmZU6gXee53m+maPRVtGqNoRG24AHJYgJQRsUXjARjI4gfuf5ROc6MoYejhc4sQxR0MYBAQ
2iijXrlyN3+4DPW47x12xL00dsm3MX6OsGG75Di9ydb7mm2K+B1pLRTHYb0fgjky+eUdwc7FymGL
AKzPZKQOgC2XUMbkeJws8K/fWNwbUNiwZD7VD5QpVonzsrqQGP1eid4+X2ndhvDCyWyLZMt5JQHB
jMEZRDSB7mQgSLP8jxgzWKIJ+PlwM+M6vuORCVFKDX8Wb6Mm1/p36AJjNfgs/1e/n+g+dcTu4sKx
JUjZetTo2EUIUTRgATUwJ3onfVCTLKgMiCJhbRX2uX9vi2+bnodf91ZfQPttXLaOq04Zt+/AS9R2
jeq41DoOTcS63AEZht0Cr9T3HohT+vTVPsLHfDy/bLkMLGMhrvI3v7i+9KuXOLThJbul6L3oKVhg
kWDC6QLv1zR4aFsqSD5URSEYwDLWIbI01W+VxtUh2jwa5l2JDfQd+9w7CED3WVtl/ahoqd4V7u8b
O0Q1lF+eMDY9lB50GumTU/1RBxz/5KyGreBc1uYVtwPdGKd5lYBuorI1TdLn/y3tVL2jX5wM0Sfi
Pa1lohZi2PtoR2N1/sYHjahUls1VtbPkboa/DYIOgH6nlORD/5v1OziXZiDSf4xxRloL0EwK+f6J
p9OMvGV5QX+EB3sqUEAdX1mp34DSv/4PloeMHE0swDysQ09a/bUM2xS+UqFqREemAiUTDT4Wz970
2r5t2QgamfGEJtjr5eKTzjw3zTWfTjiY2ZFjs5y/GD0jGj9EomkHQuO5F1LN2qmdUpT2WlkNOEyt
vpNMwegm+K9Y3YZbETMe+/4NWz4/bHSBhJ3r1qgqHipjwKvzg6q0nuKWyoRYnGdkZfHb53bih/Cz
UhhVZzVH5jQPnZpe6IBlSWB5b1E+tmtVQFyON5rI6L2enBWp92XFj1+oSEGGUW13TB/dfXFB7bH5
kMMd9u4S/infdFqPaEnprfaRxIlWkX7pt/jD6OhSVruQ7Bwznh1LfY2/cjt4YmDXtxCvcO3LcBVo
7RJy8zlEyp3iT50dy20usrwwfzCmMSaDTFYxTX+ActRQlUAHFH2GprQSTKIEMRhQQ/UASgqgJgQe
DvBZdN3dmVoEEbP3fhL1yzb9RjCcUfR2l5cqJV1wXadOf7g0Fyh2CHYwB5wuT9QbjiXXLqZa9H1t
nU6ahetljX5CfFQyljIb64eF7fsYs9HWhWgHPUok0TYRNmB4dWRZY8Ptfturw+g3baaI2HyVUnki
9Hjb8CqAUrthlCo97LHISvKzDqaXY3vGaPI1xltSdm8rKbLrfQzZ4YCNb87qlav8borG5BYe64qi
SPGlfkLBNHn6j5MQybCXNb208M+cHpmYfucy3/mAuHu8oC3wtrNRYWJSO1fe9RVcBxM8hN6La/Ao
eJsfQQv6U8HTE3jqenJnqgcsbwHaSCIlif7REckQDrUYj/pLrP7zSlLRwm2gduxd4q53OQJSUmfm
aclGA6wWzn+5Do3Z45b5t1EdCpvXatiYooOvNLa52czB5sK+d/cwO5geL/k1vqdWWmCZH1c3m3Gy
/oA9yzTVYVkdnHNn7jxMkQfzuVXBGPCsajhg/tJ3/o82sCvT9qJOvVZeU4Zw4QXH6xtUPZnsG2ih
xwRfJ/Voszcik1/Gajs1QPdu3t4sQjVYXxQkKy3WdAdT9VHVYFFT90sjPTdGe7c67XBFX/HuFJd6
Ia09cT9cwBitJL3TkqDnmphw56aRduPIU2OR32fNTisBFgcEw0RiGESvwhp6YU8M14vs8mETctZd
XzmeATDRqVVq4Uut1c86xapq5QDBjrY3Laxgr0C9+/L/Bxiwb/Som2qx576cBvGB+QtFDkjfToRp
emEWXwOKqOjoVLfOCA8093gv6lbt2ETWrdsaM6owX1FJo/NZK5CteSHBpfg9zQLdm9XIFfA+ll1A
SOfoTGIPmyw/4Ae83jQw593XHG2Vi1pE46myzds7BAaTGCETHWWc5rKRT+YGQ1xX+VyPluvXFnaG
c9eyuDRppuJ0wrKp0lkkxQP2a3/Beo7PwgGO28G9QxjL8/u3O5xfVIsfK/N0MI+81BQCIbWKRgRY
hhacHEZbYopakIdIzQPyHhgKyqvO0OVeaNgCuei7lT6oa3q/mmBRoYhMe8kHa7v2+bq/WlwD6lX2
V+RCL2C0qt8HYmNtS57F9UR51d/3fHWVItBncJpl4FTV1RC9ZDJh8bQyWt8styjXlvtG1h9Wx4uA
Gi/DLYb/+63E8PHKNAgq2Af8PcgbjalP57rzEvFzpUef9rFSRjDt/r586Oi+eUH4Mu88Jtou0hIZ
5+m5OmVlPo1s8bP02Pi5zaC9rhySp+utukAovsBFH5CF5kOGK+mA5E11yrrfST3BmFgQWcU4NHIT
gkLkfdGhcrgaL7YNUYDU/PmBUz7T34VE6y2dOk5K5y+9Du3Wm12qqo2NTwhzSW+pEuDweTwFI/bm
CSVplUEvzxhsI1Ae0rwjtU8foQqDi5GxhiZZp+08KJdgxW1pLFiZDzR5CZ2gdBLVVO4nOyJm+dr/
BzSeMwLipl+218UVtMuWQCEhnHsdIFnnGimEDwG4yqriigeqpOMpEqcZhE5lkTvIXa/D8RsPRsSY
yW/lBEsstPgNcDlfQ6d2QVhFsz4FTOM86GqkTnm3u5pbuX99OMmbUQwj36+N51dVwcOcOQ2w1Q7c
UPJ6tRHlVNZHL3WQrrvOfid4oKW2krrHBCOQDzI85X0CIqUFBxGPz8MTk/tG/qym2q014Wg62npG
6od2YjBFn2Nvb4EhEGQ7zMRvYs5ny+YLOpTwo+6NadJ9UfzCvvWfKMKLNhzWib/OiV0/4t/a3H63
OehcXid5Y7U4X39Nlefj6wezZ9HEUQOYXXilUbMrcNZTSnonbSoBMn1MwcBZdPNeItDTho4XUtrC
OhrDextI6XdXbX4Yww76IT1pdczERLoebp1JPBe+Opewuiu/9m4vs6QJFG0HW+JSBl0qkSjj6Wz1
veRs/ish2IEaj7waUOw8WumlUKh1W3QCPI8/cmBXCejeJtjfuYhSVfeh7ZrU3bPjHkMLxpjm7yYi
W/nKTY1AcBtFLzt65v+kFw7AsrZ33bTxRlduDOwYL9E71trLtkMY1XP9ViXcxdKgeTErfiD5sWk4
L+cvYhMOj0hdzgTf4lzyh9DzKo7NheXy8xjBkh00jxxD0E15ZqTk3tm8Kzs/Kh0PixVQt5fpzcB5
P3hcmAOYebopXjwTm9UMY8q5alqzfqPVx5aDo/fug8U276VoQBNRiQLP76QlfzHFBhbmYOg9booa
vusNnQI8PQLRWJkiFugN9uiNza5DJqGyw9Lc7vWMxTOTxJx83xM5/C9RjMO8T/I6ovbanbzAhMWA
iluAlEMaCwzwDTgITcZguRPgkGmQX1wB9ukFXYPZyooadE+ijzb1J2AJ1PRf9hl/UKRnZixpwck3
ppeb1BzxGbjqKYmmtVoGyKOOB8KdHCx8hQb3dhsTwVTMNSASOZE6cjmYMMo5fxkXKOkzrjzlyogm
WbDfEIHUHcAAKxu1wAtG1AMtzPAr6/Ih52l9Q6NlshP8vnKUL3OUliOyVfSKWu28n7oj48Mxy+4w
tjHz5TDby+HzcJm7la1hicdtKimU+vpOK/hmuAp3NQIsV49Z9Ex8hMIDdC6dXXsViAL0suPu3uzX
/oEwiSOcAscBvgtnTZqbpzcSm5KeEBWZeLfb/cp527MDSMWOPTRYEdUF/nBAdLFonmUaL8IFlPT0
KHggd7j6eRsxGOl8So835wnoW0XGdXUmk9ZYZTeUCKlcE1f//muRVkNeznmDzhkAFpSET2qDqhPR
Oq5LAfZyTm1fteAPzQ6NxB+G6hgr9jGspmA5MOGk4yWPJdNv8jTsoaFHW3HUS4fny44vxQwMbpWL
Dy6vB9upgp5f/Ji4XUjhROxTbkttal9TasKws0YLqfIfBJQhLS9da5jR6feIi9B2ERUwN3hKXc8y
w1pC7FbLT6/UomZ68KyE73HkVhvkG7FbBVTAfwt0w4JN96FcJwlqunWkYgdhjjukJWgZiNKj+DlX
5HVkI1z18eaxCGWYvP/cTs4yLMZpWU7ducMVMazFF9oIhmNit0AR+jCHU/rO08apE884P3zhZzWM
WaDe9Kxqt6oquDHH9CP9XwoXcg+nORHHXQNCkpu3UpKKaJ2GK8Ym/HY0mfnObvgywpyFvDhJgPGE
mBpaOSmBNc8OfMxCDyerL0vNUZeAnBzZSOFsHtBPjRWSL56OLqOwaWZHAj2+xK+NqS33/eZmmXxY
di3gkaX2AUAuSHbi2NXCTJ3NH9CdRQ7l/wDg4avmtlnHwsnpnd9MjGAsYaRE7Q5X3BuGTkyYebka
pegNj3WXVk/8nntipUWDm4u/DWDmlOqbPepkWKM8wVMhsjQQbudKLQ0opwkILFD9Qo38d7/AubI1
w6WgQM8zF6P78+K+NnBXsUNVGF0SPCiDSpKgBGePkkfzQd3HaN2BLaVn4V8WeUVxhXPndTMVF1D/
0jV8AEO3PYSEVddjVxaLKtlbzhGEgBkkUshyl8milJNpcu1bY1xipCsxNJiS7qLKcJwqRvBC+F1z
wuTkynLCbwpzodvoh1BhaHHGWHqCzVIB5qcJONdW1Nn3WKZzUNYAWQMX7FMACDWXuXxiSXFolfId
iVU3k5x178m84yQ/9xgMuROgX7FmUfOyrlRaPD2J2AuIrQ2M2CaZ9SPQfjWuRFz43XoKKYDrjP3C
DVFnZdKv0wGxPHvDEqvjeKOt3m6alRWh8Nr0+kToxRRUqRQ+k/1WSmDNm3uWmglUdWZ+LWJnsMpz
JIbhNluO06/9yp49mVRxAsRtSvcyWAtGwSbkBhyBteyy1BsYA6l803IgIaXTBLn7V1rHd8gweT/t
WNCqQhrY9sr0kp1Ubo9ww+mmVMtjFE+ghtH19TBgJLbZ5AbLcsz0tY9xe+grQv2wKt/heI9pndL6
s9KfNdfU3F5gB3AoDCf5Le3IKaTp8iv6OeV3eCG8euOwy8Cbfnc0ut01u7UnET0ilnVFKSz/74te
wuwcy+tXIIv2xvHq2JgWEEdsrMw8CZfVTX1812iq5iKWcUTyrvo9ooaj0GsmeEcPmbamMquxShIT
Gqvv72urZDkQtFiR53DYeqNKpFVAMGAXEr5PyCpbNFSWITIdCBaKZY+0NVxQh2mUrt8WlgU9BOzq
69sJZFzykUteRcgp5nY1oE+78qFI5pOdyEcipp7ocF+jr6CoJERNVvATRT0qvWfO87BtLyj6gYC0
2/Jwf4S30phvr9TYcMn05qCHga3cd2fBj06wIgLt3Mwkw2guvCyq7Gz4TF222EkhI4pCiaLc83AX
e3hcYuOWPvZM8ulGFi/dpB+nV8FSHo4IS3hUZSLSZeXERhUwxSmU8rrtFAsZIx0ofpRrSmaFOxgP
ncCPsJ1fO07tfOEuc6ff+u2RDSctOWEQL/hQ47OkR1G9Mj+5xYnMZB7v26B2nQTV/PR3KkcZJXyk
L3hc5RqcrhKR1m7DkBehaolzI0VEX1emZ8F2xQe2S3Zq9dedlaHeMfGkPAyWwyWE9BE8iXq30m8p
66eXd7vEiovgEutJWNQyAypMpIKqrPosh/CjBsaqhdrWFAmbb0IwMg3ag0Hq6D+IopjuEIfOiMuN
v0FLtwvZL12PsindWfOeCUMmcyqfGxkcDcRL46F4cWgeQVWFgoKHMtgWoXSCvPoNOwIEpTRMfoPL
fSmMzjT+GuoAraO2fr+Ov4YeAUlQzvmV0ZGxvSonXmeRJxA9vPPwgtLpQljMmBDiWL99n09aPHbe
LjxcrgXegSWTBCVfSXM9IjjN1EnJeVwVYPuoGZ/TbK+sW5DPV0kGdhAmcc2GNHPPoLZTXKdaHxlN
4nkUKgYEd+vXsiYGnSaMHHd+jwhoHp0QsS5BexUGlb8Efh8g+GBYPOJW7FgtUKUHJg+alKxxWlts
Ec1quyZzF9St3zyr6PGnA5il1fL03b4lKIGMQCDQZOekfQbpfTvQIJYHvzVoIPYYhxMhKj/ox8hG
qa8kFl2Y7jNCSi64FpUsGmmQqK6mHl9NDFC5vUXNnLIz8oki3joXlUgJyjzpu2oSKAOBGIVVAtXF
XKoEzSTrewurmJ7g7bsfYCw6isf2CnP7BXJQKSzu0VhA3XayyN4XO2neL5yChlCgY6KIKCqEx/Z+
o/j9w5tsZjW0YQDlUO2seaSf6Num1z8StP90y37WObhbWDiCtxAVjztezu4faNoAyXW9gUnhz1Tu
Uqp2Ss2e5auUm/IJKk2jCKihhlXsagctFJJZEi1TOHJVEFyWTuxCLZ00THyXT0cltSI7py7XKMOn
QBa+1AoPThW8ZNbK+ngivJcZxGwmLeOw0Em7ydWOjKh1GCZejeEbH9qhUeKbInGi23wZCQRzP+nu
xbRNwc6UuuAxsMUTayf9AWw/5fqgg+OdTDZ1jiuxJVsflKEdoU7VId8yJFvp542gWTf2VflwidIm
0+8jdGGKStaWqGYnc+k7YEAuHMDOM9n46lxsewLaVGosQusk7+Q5o+a8zM5ph2CgyeQo+Y37wtNv
15F7Ub+zfLMZrUugnab32ovVChk+zL384JQEgJcfVil0PKbqqxpqo4wOXY9jmCFJtcIh4XDfjNKO
+93c6MMYzNugXiJCVv4pISeuODO/gCK/TwzdDUU+1lTEGMnXJ5g6f8WBYN0hK/Llj3juSe4LcFcV
Z/Y34A5cL/GF57ZD0w3pdyKnjfWV+al/ljclLtzLgtcdAZthggxR/9hG2PzCU++vUGWCbc6yXQT3
9QTayTranwofQoJh0dxE0QLD8fDpL8wAaaaOydWMyfFY5uX8v5Un0Q/yaw59Xl7YZr16RX7Kraiw
Xvbt/N3WNGdG9FaDsYtf0sYEufJ1W42wGrKwkh5ypKDLDH8iXCTtGjrn6lbLGjgHf+v2iXSTgZdO
uIXX3yHwVFx1qlNOvZngYjUq7U2d1ZE207FKflMW0RXYjGXhhfOLvMuhRG/5lZm6E+XbQG09bUvc
VrVSK0/xE06IXfs2IcQtvWTDgq36k3psp5glA0mXmCb1U6siTvXcBY1L56CGSfpTK7TRf3aUTOXp
mq4SDTL1/P3exj82+kTMbsyv9tWDDimLpnNkWgPPBj5Tt4kgQwKtUcSKWOewZLR4OoNWbKwm3Dga
xsC7HBtiz6GXfd5N//jQ6PxTnjTi4vKwxR7zGBlWQqczfbhkCqfylsppTEWcnjHS6cr+ZP4ynuL+
S4fmbTWv5DkWRFAIf4tcvu25xKf4i4x/Xf3cJViHuuXNxvXPA7gtM2N94ZsbY5JWa+V5IvVxUr+f
x1f9g2YTIB36c2s2cj8nXlPZy3xvTMR/FE7RVM37vWWYUh4lg/GQHbnOOf9BILymQZorFIqeLKqB
aASbKXmzggv5YTVVcr1YwUoc0DgkTc+83fRytB/iQICNQcU6Qna30JHu5iALfPSYvz/oQogu3gkE
t5jQqGiibGEDd2fzeT40V+lDTnNKRWi1KHLLvyMGOyRaPtwZlc2lIXJRa2Gy976/PLjkJP/S3vTJ
tIQvd4YYj4QB/EkxzaI0gXdN28EE9V3jiyXQC5ktbVjBv6PKfFMhxh2yUkYmyJfgfZ3TfK74TjuF
aMXMIfJa6KVALujUf75YYLIrbccWRjdKsSyoatbVuikq08w2KGQf5k3ZOg505vmyUz5Zr2C8u+yu
Vocz0+6yN0dxsmBiikPczyynHGeOByxzrcKYArGqFu0VvK+0YtBJ+c0Mub+7gVk8/iMtHnahkjS3
GF3wBcWx9yfzY+fFZeQNzT1TEhDe7MtdF6y/V7a7NN6AYaqZmRZBUttg+Ussubt6yGBRMOH3hi9e
Q/R1rkcks+eB09YVVXydt9TpPqzTRJnpwzV5Ct5rQ4wZpgNcLGuGL54tYkGOlw3rgi7uOFKT1cOe
wYz4sdMrFzJaX7UNzcIhvtQ9bZKeOeC7fP0QsViRQvXJAP3MNAPUrKQiraoy1WBU5nDNLSgaGAvn
xW4YtJRij9Bittaw3/0Ox4vH2kJ6PMkPEh9KRQrOfXOu73aUpwK9G8phzF+XgnwmoTYFt7VYtGNx
HoJYkwhE6SxNKaB9VUx0Y95KasjHlbiGAjBmHUoBVwt/bQ+7yveajIPMSZpfiu/pFvmsEw6Cotwt
pibKlZ849b9/56MGe74yuNOCATcgKV9UZ4Y5op/zSG/HgvHOzDs4FXuLUWi9PNKXfy2f8zwChRP1
FXBK5syPQw54y/tupap/siViBfAVJFUf1avR6Bdk5PAqRyN4tcMIASkagg8ZncKxxSWdxlCWj7ta
QCbRBZoiw17bwhWoivDSuNBS7lKiA0gAdCuSHUNXoJife1WDyUUnmP854KQcdzvglEAKQYqqsYRJ
SQPBzTaKWyxlekX3r6nxGObQbM3CDSz2JI35Yya3myklOwi1wpEqrXadBvd1/VAsxQGpOlLMuUSb
Z215dUsEWxAL5kpKCV2mV/GpwdnBzYKBFCh/4Etm28d51Qv1ZTA40efpFCHg75ZT1mCB/cucSt4I
7v7O7j73IqH27xQ/jBjiPdThfa+9iZOytvrFEmLyl3nQtgTrLC9PZ2pDaJ3DveGr7GqH8QyhdRxE
kAqejB+tqKF+MGIT+cJhc03srjuTFggNFXnl9gvuRF/KcGtkJMm5fmYP6FesOQ2oIYqtWDsKTp2b
0QvdKL499f8HZ/9e6jrGklx2R9rn5lF2gEbgrzLvVzAA7Mxk/F8y7ORMxp36WduiGRvGj4zYsImz
rXvPlV0WPtE4RGHORk8kkTUp4qEmt4tCiLmor+dn/OXz71CMioO/fj+YsM/CCnesBOBJgsxnIuxQ
iyYPk68wqHPZpz69BsyGPgf1CyONsE2wUhPjE5pS3AXuHFN5IvsXNqlxVh2dniCbRwpSDqjJtdiD
Lh7n4i9E7sdifOvsMw/k9nPOPo/udr52y28/Tr9I1mswFi3DLV9jqwxYB4WH/geNpXEQUQQZod5E
KE55D2rPT2/VnfX1oWlu6ZEga4LGxLVS/NHr8FsYKYKB72tC2FCUGI0ewgloUh/66gZ/zmKdPyRV
3dLh1c9/q9x8INrIJcMntkzX0xBZCicDWE3j0YJogTmGXg+2+Olkb3on8TaY9xkuo//NIwd0TK2l
Ne9U4Q0KrxRapBvRRmIgREyXbVYAiTcYjQOjdt3eBgTifea4zkkJwXny5R4KLGPDSdJS8yzc8sjT
ouJCjY0m7Hz074nbyLeLyH/pfhVYS/V+QaF6DRHmOPAZTLjjHr3zTwete4nK3aBK1D0s2AP2ZHH/
oI0FN1+gOd+nOXGEnymua3kOTteQwae47rAWFMPOqiRVcbwxulux8XXvfIB3Lt5txBGxbUKQxuz6
y/I3o67p15ZDxjtPZ9EwD7UKmOR+/G9iESPRAcBQ6Sndm1y3V6WnV4mE3NBsZs7X2TM5YN2UThjs
jJoXLkqLh8VQ2ZQ2UvQ6NXjP6AMCMyK+/py4NwfFiU1sDoI2MXyc9i354W8ithmpin3cOv5g0uuv
PmiVYxaMf7HpDR6CbExtp/KHNHCkbN/gPxeFQNEgU5y9c0rUihcc7SCnx3dGgVw13ldPVlblpWHQ
AE+KaMij/NqvjdrUM2IKjaNiHnzo+pwhZDnm5LTR6E4DXXKUBP55qtZyQKoodrRV081lzXTCm71L
+yFJ2mRbnp5HY2SATfwW97wd7kPV8oWCkNII1/L1uh+FhxnHL38l0ycbgZ9K1yRLzz0NQHxzQ7j/
hQ85/YOD0Cvn7jAnJHWHwDAll8I9PSF6s1F1gIhqAR1vpr9aj5kbpz5va6MdXj9uFuCZbj8Te6t8
BycWpPOWx0/CH0fLydhz/31QDjlpVODYtDW4LHKZVvbGwVJHVbvNFlCZlMN8TOVyDKvQOzALuJ6S
NfbVSoBOhwM53KRdRBk5SG4wbAY0RmVRoam8xQcmCsavPIQKFrNlBcwMXGLjhEXvPtXPa4v0sIWc
zFycJ+5Munwo6ikhl+S4lkH0bz/ijVObivSufEiAA+cxJToEpSG2k9e8CGggfAuiCKyWnz9pmLSt
wr5T5LnQu+B0ValxPbKUwavvNqKYR9d2mGzFgu+m44ypES3acwtcw4Xzb3TA6np/iarBqBGfM3aa
v1/mykMQzb7NF3VUH3fyB8+6JiM4ju4MpgTcc/kcqCmRrzcsIhkdwndAb1jfdPosIYLp6AYA/fZV
FIpV97oGyt+D3s5fDUGZNRQ7ySvbJwDLHExvacjISqZC7m5vP2Tq/jt6wqmFMSSN7Fl0mhd7n15e
D/fMk2Xu5gYo0mYbNIBCkD5TAByWEo3jMakXCFgwe3/F1G3g0D2JUA0QmvRB7FVe9E/m50kZWri+
9ZqeD4hlEjZ+8lt9Si5+n9SDcmyRR3KHA6mNpk5SOVvcrpRXztwU04hsYm/4WKWBHKoe6j9iYAFN
Yjhth+hr5QqNFyl2SkFjXnER4f5nhhdKgQlQNIC7rTT37q4ysZMqtrR8yx4R8kNRajwDCK/NnljP
G400fxJrgFkLlvYh/CHhnkUTgwRTSec5+tnADSPRcTNRJJ0KjoI8crm9IgaJt+G1zhtshdufadr8
kZXdE6oRAhYqio3JnZc6N2sS1ZVzLE35e13DLeK0iFKSS/olE2/XfxlYvKRKOPq45UtjWz34oG5F
F5YagPd43eRh4j4Capun05z43ChOzLiP/VxDt1PJIWmO+96f4jkX2lJUVDGZYi0323B9CwTygQK/
YlcscmWd5sYXc4Jfl43QSKCeS86jHQm45uSIrSqUn/vDfWOhECa+cqPp5Y8X3CPA4KZZeMop/olp
vqxYk7SR2ZntZ8HjhiZ1K6AKdhbjqjztkUdEG1xcmY/6mjj7E8KFik2TQRFT6SLjOQM3ior1yMXu
4mRMjgEgB5+KO7ewZ8IfffszN3MdWn/z4YnyrLpMnZJ25JNEI8p68Lfwq45A2y2RcAEg+llQe9wH
ID1KemZlpDhfL0mF/eF/bsRSUDgCFuILsAteofgGa0idHT4zjvA9ViAR9yTPALjhXKEu3Dbhge6n
WyBXA6eD8m5RZ+WFKrN6NFndwSSrEHO2Pixp/zzodxf9lN8NhfJU7Kyc5s+iOr0HnRP0asQAVof9
9jlT44Rs+VVpCXuz+gf1zzjXexAVO9U8bJ5EB9Iiovy3fbLmIu9UbXKTQGnyWNLDwprOIAwfu2ra
9Mxh1vaKGclKdHgrs4ArpKT/lK2l92RRUdd0tI68uDwc4IiRDCjN6SkHuMiDR4ngskGml1h3Ebkc
6NA1S0sa6I8Iiyp0R2PQYlloI66CV3LqEeHQ4vjWACdHc/UR79jH6F0JNfE0gahhlLh/l1geckgZ
Sa8HWL/+LdFrtLnKireHUnPzy90F6OAt1hcV2fuhI36VxsEejoBQwiqfZOKlLFt+Yao+TYBBPsGq
vXTFWBYR3E34Dxmx+XX6+qDXQUp00BfWwosc6xxuDrC+qrj/trRRSfuP0TZYvvo9S+tJaMqSSN2e
A0HhA6T9yaYyMROMb/fvz3vkTpJaXTcA6Za1BOyNX+pq5UrLBgekRTYxI+Waa5FaEW8h82c26JRL
UsrZvoMzUgdNAlHOMHM08Qq2EV8jAwqkptJ1LCWYfZv+Uo8G2oW3FQpg6V8iAX8W71y1CH6ZXR91
9pjae+j4L5q/BAnNKdfUM9IqXEhpZX5FCAcGtxv5hmX/zwE3HmA1CHmpCquqbtmKi9V9UGSjAh8C
7sj78ssg7JOZvWxcJE564lFm2fIPAba9awfMbgWzeTR5UL/abzkm0RhEj/GOcMV7+rIPrO5SnYPx
JlP4iQSNHSn+LNs5vmF/9yZ2ntOD1ng0Ofm/FsMDQ+XGYKJIb9WBrP3cuyExQGjASahv3jcpBSKf
P8fMlFCEkTjGngv2WvDqmvkZnk2P4T/6+OVSFClkNtu3LnIReKlOOa5pBQHBqqia51bSBSAj9Wu3
VphNP62S6+QXnwLgrpb0AJizjn3NJmhu4cmmXii0O4ma1ppjtZMRLLf5V3jMQhniv0f/lzQqkw1W
jbdyCQYvWPVPl97PQY0L0x+88oug2JUDczzuWXE/iIqOgltRvW5FHhIhG7DwC9ykfLh9RXQ84KvN
4Az39s9oAQQJIOrEAW4xtPBT4dVFmV0Wq3OVBDeLvmjk47aGdDFpdpQgCAOsDTjs/MC3YcWzuGW8
AkzlSxufHf/tXqV7twAP4bmzCq1aNum0L/UfyAAJnFWWrWL7Pno9O7q9Ms/Nw9/R3Nfn1kuxLv6t
MpmVAVCYDVHn8sSoa79YYEOVAChuoyS/h35IkI59nwqkKlZqqTkZauxTbsMHpPKhR3lNtjdDnXGa
VRx1KlfYjyw9o+L6+O2Sy9zSY/jw1dyRRkUea8xh8ymOTCxQFgGLfBuTO1VYSP88aLw7JDexM8K2
v3HBYG7X8qjk40a37GXLlKE606BX0kiEGueGUHcgYNp8+5m5S/eJHh7yI7yTV5a0bR6PHL5qZJ3v
36WWDzNxvg1v2DIvFkfaGvPnlMCUsscBJefP81GbcPW3J0zHGXVYOdnrRQMg+Slvip2xhv15tEDN
ABD/roj/LqWGLwTURKlaC2dcNVw1gxv7cIgidgkuNit8iUYAk1mLykZQbVR0wLMWT/VhlrlI/LCD
kAiIdNJiSM3Y+fjKJj+fDJ/QNLn2Yt6/toZ4t+WqGzN9fdo1HhP3YTarCZlFBR+zxr/AVAGvE5IH
EL/7XItHQ2xWKd9UdfUQnhOUxgxu2tVKY2Riu6f/EjKafQATg22K4VE+DdZZpMuR1VBxK5PtAf+Q
puIwxL8AoYE/1e+LZO1L4SqntweuGyUqzGlYiCc9UHAOAngJHH48zqhIoGIo8np3f+wMw1yultpi
EXZGss2fus7zCKcUOT6vHDy6WX2aHr9ej4QayAOVQ2W/f2BweUfWZCpsgB7a9wjaYB0BtjxD9tfz
mEGlsaWE4/OAzlZun3rf4+a3bq9uZateayxrrdOy7Bkv/yIAXr69ynUBM2BvkkUl36MKpVnzW3op
Nnl8F2l06tZhp/AQTw9PJc3KqHx0hCqDbpb0i6Gnvcfb6Im+35+T3R3OxUpjT1H2J1blQ81gT+0U
5tOXuRJR2qpcNkIjH4hpDGRd90zsdpcesjGzwK+bT9spQCglzBzbitfJQtHL2VsJRYDzoVIWiLKp
2JJADtke+U9xJnug4/MoUZnsrS+PDowhAJhdpKBSXIJUM1nCUs/GCoRFiywD3dYvdSKaNtki1A/A
h7TWSaxZA+8c5du1848P9Eu7TAsYtdZMVnBbO5oA18ZvHX6Z+v1sfyRRpinRja2k0Ebcq7jht8PN
7VGMh6Zl19+ORtY6iRnZJDkJjMC+6Zn+WRHfWtZQx+ztBeWs8rOmpw4u6/x2KXN0PP1yZMCCflT4
uGCRhHZKU2vdkkOhewv4Y8mqptN+R5Hq5ooAmpbpBkjGiTd0Y9TBJBG+tN/w6VSWndR/AVrU7yhZ
Gcy9CnMT5dutQUVvVTFfRuJT7jcPI5AkGnOpAtLDRFcba1uU6H8h6b9GL23ViQ4kliCKS/7cStyd
fa5W+Xi32WM2qGq66tlzCnGRCT2Lp+o/qF3ob2NmxjH0GB2FJG4xiOkFO6IcE+U/c6XrAnCVXBx7
lBpmVHZigy2aCkfz+MYc6yI/0FOWRLNgizdgVF/quk4OAq5WD7yI5DCwQJKLKQACaNYx0qRS1nw6
NbguB1NBs/RojvP0L/Xo9Ci2ncYLWsn9LTWAH7+QUNrv16CFa/loYDB1yV8hWURksyZ0esSCAiKy
GY6HLuYR5/6+4qHQA27w+ckfUzHbH+ae55ibVaEl5/ZaJXDeCdJyF3qHXFFyWvNREwoqH11Q3QdZ
G3GJh3vqeJB9A7esnf92EfbdZfXvUc5cnBdAoZBGB7xg7vKL/mHiZIG4zevaTAYZAw4mQ9pLGPIL
bk1yY20MAUJrBW49Mni0mDnGj7JaTkNQBkyE7CfSNvZdRYSAuhCJTYg1Q1CDRn8ATFZoBDzk74cc
RAHd02a/O+mIrV3gwBT8PnbdvJkguFqSxPsyY0fVJ90cFrmj3YZxIdNx5m7PFzjKYpfT9mMe4TEj
epHwYRYXAXbFkaoW8tEBTk7AZAURlBTxjh2XhwJ83gvErViwMoUny2t1AaTyki1NdVYEpLB4DTk/
iZPtj4uO5GRnKrbUm+KnOUltrM3sZ6wo1YQPVp+CozWGfJjcISxydVV8DbmjDlpHSba6Oc+fcFxZ
yYYzlpIpENJkDImNyrwMeqUruhkm/6nxFkFuEgPZCf+g6n5ke24ncJrEqSPQnZJiCD+T/3Vprkj6
j+W7/AdeWfi71KWWUq+BmWSwEKvdGJYRypafDYhteZ/hMGUO2wD5EhynWlYpF/aPxGX8rr/3qTO1
s7dENUkn1EHBdH/AIGACylu4Pp8Uay8p6T5RPRZXVRUYy9o9pSQpnhpz1jFV6Glsa3x+Wz2SsXqv
QSeEHEdxz1lqJeVZlpEfAwxwHsVrwIj6ChtIEeI3/xtcK+EgKYY6BWLf2q8ZPtqg6xDukDZkWavy
ahYp7JUEbEmUDNMrk8RfwHVjcEdQ1/82bey/TVlrAvp9dgrGDaxgUPdmlOmJD2AhNdPALmsCb+ya
x30sbwKrcOI/aROyziGYInWwVON/9+MDYPnFhnj0P2FFDPDNLXBk8jc9oUbEd21bdyV6rN+ssD3f
PWT9+rJt1iJyGzhyH8zElxKICrQHAohYjFK+zDtf9OfEyW2KqC5D4S86K9UQcwXKji32DsIc//JO
ANwo3tr+Qn7OHGe0WznQlRiXmW771ks5N6Qfyvb06gXj0FM6zOHWOp9jOiA0ntdRQMg/XxLXSxjc
hrS/yXA8DvmoQnzvr/oPqcUracQ5fivV/oKHF94g0zgObzAQy91chr8GVyUvQyA8GCVawlolRjgI
tPsItSd68Z3+9ArK8+dlowafs6cZDhC9vP/V4YeYqSihXRTvH4IpsHI3tuoeAdqTHueEm/3OVZC+
vVtJDxCb3iT0vftQIYR4iDcqTBng2K3JFHcWF54Ifm/4m/NG5CcmbnMJAAuF6U6cLKaR6TSSPIL3
0yWkLe0VxoIdtH5PrOTcD9FO5YbGXq1Ifk55VWKYayeo4XZQDSlzK+aLYjZ7WgMalQCAZPQndf7M
rqyg0EeopEXEC7IWHgzVfvQAfVcAU+7RVCffNHdUAsHJDacqQs5qW67N62HDB2mQz8hOtYpmwg4j
ioU7vHTwONk2aXIsyRUqf/cNtGzvEEvNeH0eQ8kuT8F+BwX5D5wXn3vaRj2Zbkxl9Zn2Dhqlwhpq
wTIBmOQyaG8eMxvbWGc6K1LEbHCauQGFwpMAZ7IZbiYz5JhzBNzPZEE7CeEUZcYAvw/062uwF/Fp
UpSSsoq0FpIQjpvEy54KUbgOQ3K7/eq58wLr6nZTphkzQ1B+R3fLoA1anF4OIXKi2bONq4UA6XAo
WXY6OkR97snwjovNbyRcsFWhIMTediqWvy+8E0OdQvbXziH2tSneVUOb2xtmYVnBRgk7qD1Pnygw
U2V0dsgdLUXpD99ysIYb4nyhVo8YzNGd7ejW3c7oBMFobc6GUdYvC1ZJuNqeyUTao65Vgt2rfuLK
8bwccLKkItQboNdVLHAItRtW4IP3O4BIC5E3bMqFfg5l6u/zVSxsPyokFumdzlHQEVb7QYauZsNV
fC5d71Lud7HjpfJhoULzp9E6dbMR26I7f6j6lvnKtlLTRy0HwrDMwJqJYHhNcpVnpchuRv0x7Tse
fZpTDO5epj5yXkJsR79jVZQNFkHu1xfGLEg6za0e77q00Od3PampnPac6UbN2TYk9P+W3o/mmkeq
R1Q1GwLQUf9j/HqK8bDLvhCugr3xgLd/KGXbbUwE8/sq0bou2gjaPkcHZM2RWEwVvqYmZgwKGR0j
O9AjbB74uVtMCg/ew/oPDOiT05HmEu7kB00OzoS1xtycCShQmBRtVrSDkvHmJspY4LaN/K0rojBm
xjEMzouSHEWnFxHlwHcUlmgo5IRNcVUUug85OtdM5zUgRU/n/bqRBfYW2E6rP5nsNmyW+abs3vJ/
rONlM71dyL0GE8VShXfXoKReo9INaoT1WcqMu430ojj3LKK+N+ZUpRxf59HR/wWEvqoyGo/iCDuZ
7QFOpgecH7x1yOr7UAvrS6d/ANU8LAW+HcqhMAj9P0yxK7SpHEUV6dm3LlRoqkzZAIfqb2mdWw1N
kGSMNTaw1enBSVRsE29w66xcNdoBLzL0pe2q6B876GOPsKkR+OJUvJNt+1OBYJ76yrVNRme8EVNL
czEWoWj/eghP0bAlYiSlr4gOJ4mK8MQGrrhuyoWclLe2Ej6BqtMsJbx8rCVr69855P0If8jblvDw
15rgXBvxVcEYj2416bZXMNMHPo2ulZwK0ybPgI2qqT33CT9ka++1EguYeI8VW26NtW7KmohgGdOV
fj9gPxrxxu8RHCERgQ9ZB4lGH7gXX/KuS14EbeEKAsYMVYfPGupNgNUFwJuOtRM0Opv2gYg9CHNM
vSfNzA553K3Tlhr4Ph+L8DLAVD2UEmJ0ui2ukLDP/9bu/NT/C7AAzNDpeFQ6uEp3DexbjL1bFNCz
NsBECmhrVxxTtv1YbEPuZR2lYzoMfGpbjKvaGXbAC/13Jl5EFqFdsNPhMVChIT5vMIKupVndl6Sn
F6/onq6n+yxmKuDS1aTpOjWcYWc+090vScXb0hELqgBFBZ3MpR4ObnyrrsiiRg7a0n6dlVKA3ruT
zUOGGrKXlsdRUOLSmHYGElVJ2HLDPaL1YiHvMNlBB3U3zqlkJbA9HkWc/5f36XezQO0toK7ewkJ5
IFgqrYdLFecz1bwYRJHUd/eyzqei8Zb076/7g1Wm9E4/HsYODodXMznM/4J/2zL4MfRRMyHaeILo
XsVWWoE5PTam+pr3AG+bC9vvpIyEHqdLqmOqaQAELEOjA+xS/IOjPL6I+Zxd9i1Vb61DQhXkAZh5
W9CDl6VkmUwWVzHZ4HiFy64LC4aZdXpqQPBN7pcEk+71GyJWQW1HwITjsLzusSRK7CLGmg7MPuDw
qynbbJ7N87rzuIadIq8QdBb1p7IIt6ONiFZIhTOOm7moT3RNtRUKhErBnPA02OtJeOdl9IEK1XJo
H9mE2RxNpuZslkKn9PH2KQyedHNa6wfJ2zkKfpjFTGKr9c9wSABwMze5RDbOUgJBjiRAXl6z3+Qk
b3ZZ4iMXWGdWrQJI8k4dMoMxaIa/ktpGh1bgWRiKj4oKtzrmmrK/+4P2NULFBHC5X8om/44w92v/
CbopIQpqPIRSsNigHdvKi81BkoRPW+jlCtTyrLeAOVOxSjIXDV4Hm+Kdm2esSA84jBjvGCgzIOJU
NSPVo8xoI2b+9Bxi+dF6A5EGGkhf+YGDPdAvEJ5j3/MrLkXFYi+R35ksrLqHBvzS/QLavrrCoqMr
8yp3lvAWkrPLuudhx+PxwmI6C2YNLXxxhCjvHgqgZikyLcxaUGdMajKa0GTkvUTwIbolj0hoJXY4
BaeAo8QWwculwUb9zNrsxc8el1fQk/Z1qNVaGvBDc2dxvXesCQ5Xu1YwGc5JFqwgvP2/HEKxKblM
GB4ikuQ0ln8+J5MdO7qPoV4xUG7tuc4fyJtoeMNeN89WCIft7vD3bdsY5+eTf6KIW7ihAUmV6fAN
X/V+NGncxE5ODyp9pdKGMTOWC/w58icLUc2SyQxWU+MWQDvwCMDAvzeRwhNugC1NkupMf34+/ELc
ip8dCJr6PyjAlVbp15EzdSJ3H6SGx7N5ySgqCkCRj1f4LkK17aU73x7SI8o2MsDgZybalkUXvGlX
W4jC7CZXLlOwu2Wnn9uluYTtj3hDptmABz8IjLy6sLtsStuU09yyS1jtE0xRuMxy6b43wtS6VuIE
DAiQLS7UwhYsMIpKD6EfdW1LOcaXePrdNl0h4ry8wOU3tRHYsl3FPXozA8yZFnJffGW0hBIZx9/+
tDIEf3XVoLN7OPDlVHsy6yejq4oQBVG8AlJ6PHlDM738GhT1wx8ZNcXKoK+5/UcoonFkjD/sQ/yO
19BU9e0M0OOwtN4VogiW3uwMxl9MxvpAZ8c5wCQDOgYsR1en3prJmCtvSJrZGOzI2RYutI/h//Eg
ftDOSW9Kj6vEuzFYnqy40ji0POO8+/Y1XgovKG9tDGSOvPw96esJuxMvOn9Com11MK0wr5YM6N/E
sDkjEV1ysQK4KS7Yo8QSTjQPUfX21NqAXzY9l31gGVP+EHFrI9q++Kv0uCguLwsOB+816yY+Mt3B
9XCgKrl9YsLSzLsdyzduAGffz6aUTZKP5wONH2viMkZxEx8whGIErQuZhZn03pZjYU2o+fiJOz3d
QhF7WsF7dfNpu1mFJFZuB3n1g5jz3fDNmZCU7lcVLOnf4ZH6YOws0WR00g3x/epGTISZdDdehpma
G8kNuug1+xvnJ2THfBvK5H4UoFU1JZt2j7nTtEhTP5L1C7hLauScx1gI8e1opqXs676E/mfOWQHE
0Eoww+twApEkKt0j/CdPgewjFH6jNW6XyZV5fhLe4jm7kq5O+3heXIAOKrLR+TWXakiLYhqzN/lh
qram3AdJNtgxgwqRz3EHm/0ntbindmsPFl9AwZ252jjn2PZbWP4JQzgR9uFxUcs+pDrqen3jPotd
YqetOboTF8+ROmfggHqLvcvEMC9b6l0DZdJhCGjXrO8hhRimh7srLIFko5+f+snbuXLPHKxZF4o0
Wir4eg9rCUGDV940gyXlMU2wrQWYS9FZC5+YSESEvSJEi6JzSGcO/LBK5LdDJLrJGYwemYY8uZ4D
FU7XOUBJ+C9WlR1e2MfKHAFbw8I6ycjESuCYQv3/yCrBPhq3KDTDp2mcwGt54oG40hT+5FyIKh82
inMClrP9L3UZuGd1TQc2L9jVxSenZwYxDQlJ8LlnEnmAJjr8yPHdcskKoLEnIQEVkv8hqiU1+YGF
1z8MCM9WRddnubvymehiDN6fsvk62RStUwP9hfl+8m+FPhp9aaubwQ1yy/f6e4UoClioy19kGR2f
W4rjIORMpT12P0SMzKZdOkTp+HVWw6qaV5vwrwGSIfAvgNehEPOXjM3wZX9L08OWeHwy+WIP7upp
MC48mLCSilAoOmD7sP7APhNvM6T8D/X6dI1J6+hDVwLfks1DtO5CSNn6Nu594w8OgxEQDz6H0tD/
2Mghky9bbT2jINOJ+WJDmGeD3DgWjUBYoOoLYavOCNCuOmVwdQyx+31nsxpe0xqwE1cXm0v2Vb9n
xanu9sB2m8H/Hb0DCBPX94OERgYHwI46J1UXlcDt+tmi08o3wQ3wQJ94Q6Zizxj5oXT02M8vtxfy
QDMAzqx8pXEQup/z/Yz0O+OAOHvBDHqaiqM2GIMYQWD6HZwSCGUT063ODGmObuSKnChOW8GYwWQ2
5MmFEf47vf3MyALjfGTgBQi1G/wIevbY+VPbxWaDw9vv+/vzWyi7ZykwigBPUFzp8si31AIrTFiG
OuzAKvfJ5i4d/t0hZS4501o8MffFFyCvnOlmyqGMOG2tLTk3QH2LaM3jQp6l15FRXrMT1IU0TPfT
w1UC22f/K96LG4P372gIea5XVAmvlD1wYLvEw7Zp9PJGugd6M1tEolYkubkO8Jb1nE1Sk724cleI
SvBntPLSPMhIeMpXr+J6/h+juaGmXyjH9HGQ9GxlRG5sjKXY4LdNJQULtE/ezStgpvhIjWZKgaYQ
pIT/HRbKfEBnbutzweqS4Vhyh4MQWU2L5E/ugnyx0Rx4FlPyWMpFCiUhK3iYZLwKifK5FyvuEXHU
/N2PXnrUlyTeQD81zS8n4iVOCiNh5568MdBVFAZd6dHUYj3VUx+S3NvucrqhlKgeQUkqGMPYwhOA
S/R0qwKiwarrYsY3JFB+ndjLrPMFcTdj8oApja0YzA7rEnvIi8HYBJSKsKbjsPvmu6DCBz8y9D4i
Fjc6LxR2zn1AMyzlR6nRB+wg82xqcmoe8M+qzijbMSyd3s0Ffwk04BhodumIzfyHnk28qoMJObM1
kYb033TTl2NnZqU4Bur1S8HArPfwgbbr66czTQ5fNLXYYngmaK8SBlbquyrn/YpfB8Ky9UXtfFXx
usIrRnRdaJ9ksYACPZXxcD+caEYajlTA+YuyapDmf0TGzefPY5kIIxo2pJxtnLK4qLh2lc6FVhj/
2ljTT1YYdNvgjo/5jQxSkI1xDgKExUVI+3/JLtl/z6knDYugediTHswGYr/o1u+Alk42m9Fhnew7
P87Jwt+rEIIzyDOz/fc4RH9VPAVgB4jHLViYs+MdEIyMDxJxF+oft3KGJQbPmG07kUbRmfdZFQSo
YrX0t2kYaAFLCGEWL91tTIfV6RKzDdDAVokEwjB8OZd8EBCnIxQ16s4pCpWI+HJQG2w7cofT6Wtt
WIP62etGVlcwq9XpSLm/qko9JvwqSoW7HeL4zA4VMYWTIEJma53doQADVlN+USNO3n2wxmQBxEJb
w+CotKn23D6MLdVkyvCra7MWH1/tayYvAkQ32ZLTMAhAxcttKYLLlBZ9WzD74hJmo0KYTpaQsnk7
4b1jH+NFaeLEFuiKhPVxlx1I41Zw0rUndst5lSbBqhBU79zHRMKcF+xkL3i8vnwIkxHbMAhYG3LY
uvpu/bvtRZhOUQvDAAf3otAUOEbLd+R0xeugLV5moVAWOFmGBc6mtArB3Zkfav6tJ0u3yHj83KSm
RYBOu5zqGVomSzX4iL6CDDFl61nYUpjvM9c9JFM23TQbMxszeNWjLijkLeXsLw4tcRkg3qS8ELew
0uWS902c4bvU2UU6VuSQ205GRlZgMOLdiaoVwUsq1v5lM7Z/IefJWNiX1DxD6MTIZfZ2xrUH+LIR
gG4+l82PEBx9tiAD+a2HGhknab5s+5cetdDXhUr5zXWYOFbsmaBNy27Mi6h5n12fnBtvrcyjpBWs
63OClInrl+xBBShNourhx9W6tUbcwjKjEYjn5PKoOx5euf3nk/pow5+3QXKGRhFUwK2FZjDUDvtq
V/b9AI3Ucx2S7WLtZ6GmJJQE/OQth5aypc1M32BgmIhCJLhlo6mhsZWkuBaMOnaAg9KuEIKxxB4F
iEGIJ9tDoyQL5nnJ78j/PyeewhQBi4XNv54dRPr8OvufOKwvFnTNKocIll+GCVpt8vPck9ER9vyv
QqkdRMknjqIH459tMvr6jlyD5dtYqw2F54rpDNnRIfug3ALBCDVbFsNehu1DRP/20eO/GJIzrtLT
VCXq4bjvQTijypi4IFO4d6A9iR7pjEculymg1qMEnJ8VaYj6E1txTA/pNsuJ2pPZshNOhggyLs/N
X79BhQVjus0jvifwKtQGxkE6mwkkAKW+h7D6oUnRs/xk+qEuN0R5zOdtRU2iGGMHBjZRQHqXISUF
qNToPrip/wAiSEH3jvQ0AOOZFwXcWHQ8nU23p465+JycF9g8Qf1mtAeGDROOvLWJoIVDESHAO4qr
HRIpDdUDVnL93szb3+iaY4TDQRuyOgQTeAkoHid5U8FH7bgfLyoRII56ZMQnEKbRR5D19ltuUBrk
QP82Rlg4ZuYf7XYgMHdCWbUMdQWRqA4B63mlb8vzuVZceNw5wQfH+h21UW1awQYF5kIvsVm0ek+Z
kYGPnCCM21QYMV3BPipoeFBOvN34s4U13Mgr+P8bMGQ8pfspbyQ0MXXRpnF6AoA4Cbu45G7Sk/pK
J50nR8tiNAA1+eBuUTIbAGxnFrFrjfxk3St7yD4/guKy2lDzlggZiY/tg7U/RFQyF7Slfzy3lNuM
VGU5sPwvY38wKZ1yCsT1g6u+edUwzmFiexAAFQoi9AKDzaG3RlrvDMnZuex9TZrKAF5WdCH++brs
47BBT+CVVRk/9c9s0ytYb3cA1cW05CZu8xKckHMDYC2IU0hEbd40W/Z8Le8Q9xJxXj0eC6Z0bC8y
6HJfrbqT8SQKpV1Up1QQICd5PSuugGXVE/2hLuGQpgqmkQbD633j6tyvbb/x/ap6FX+UfPtCCG+g
O4JnQv5wO1bvtyVTUTDvYVNVLpXSw6PrMU2KoPUYP0itQ9ptbuGx4h/GptEK15xg3uEA5zZTu8NS
8vYk3wqeztj1d5w2sn5LiA0i7ik6t+mPkejX1GPxnfPy1rQ1u7SroJaCuqa7vWUIqojWOnt8cFPu
+CFH0oPHqpUyxhXEiYO5veQMNr97bTrNR4djU6PoDg0kBxOQuz6nqWnwNoZ3UqsdCiGxH3vLSbc0
84e0zE2klKKg9EKSCMeUtKiv7Ig23bfpU+B1HJZlWjspHQqHHfmlQhjcJAx0wJSECYcE3WjkrLt3
QYyHd59O1OqWG/3cegrpHNKx6h4yy6awvqWQKXygYHxruXh05zq7D0/qdYAXvv6hO3g+6U9Kwxct
H1kIlHBccynd5Z5/alWxmk5/Ez8EAe+fLfe64jAsFAr99yVx6Ku7zG7bqqs4GZOOhdEt//Nh+Kfo
HAlfceRfGD4/ehObBLJUZK/BcKmKaDT3KaykpE2SWxL3E6yqIGY1tTYnyOHrWtR47aXPWQ23VAIw
xS0Chu7nT+yCn9LS+ZbxSpH73u+JAl61TP7W3MBp/Cefb7Xiz/a1uInlywvrAMagpAy3gF1MLK/u
pxhNYHmXrwyBZNit4UwscXu9yr2r2EvdxnToH5ucOZ8CJmr3pEATatXiEaWPvDXmq3PQcXPNOk/c
OAfrY/rA+lUvELNhyggvpqB1d2OBy7QO1nIddoafvBn0PcRUMaPDJYpBNsmCIy4I2xBw+yTFJRZE
lgNI9iXOKTMpsEb0GafF/zSce+AlQwl+bO7XwrmIgMJ8gthcUVogKASFENLo+wXpSnW7KxQCVuIY
goiR/Mf44A/JVgwkCGr7CqJNiusEewCGr2sUCw+jJmp3Gt7h+ezgQCong0V1Rcqr6nHPnliZVfod
qw1KU7YiK6MMnZaM8kAw9ZAB7NSmRlVKrtPJ+yomS5nlgVoPv4GM2EEbggljgtPI9Qni8Drhx5Mg
cy6YmExrPL1X3C/jjasxEGsJJYRSM8Jp+XBtId9x4/4JuZMwnKuYbBBk5sYBNdOgxh9oUfDt9f4w
P49cmDrKSvyyJnbZyMqD7ptbhN8kbZDAQbTVsF4SxvoQFVpRJ06sotTRAbbQ64afLr8rORc99yy5
tiLGVIt11GI2pqnJHm1PwP2aQeMdUWrZE8jyp3SYIEE7cot/M8CrLRt9SEH4+fArpqCEbChy4Zps
lml+sJ7+YWcdOmSovBwjP4/4spQEruNDhGo9SYRWoyI7gF08ozN9NfXTUFk499jfH7OVJ1BDxdv9
R1a1bP/bVAVyM6FwD0jQdjsK86ZHvZonYWivXXJYKGcZnv4G7Wur7v+40IeYRJC8rJaTVOGnGt7C
HK3k3E7kNgA49CR3oS6IB/smKI4liveHw5FqikIeVbTEmXlh4v5avWwpDU887lK7+lQ8LgnyDRAL
xcQpTAWFm8s02XchSimmn8UYOdXVV+60E3OmGdtBi4S0alhMDIrhkkhgmNCDZyhEcoKeZ6mTfyAy
AAKbdteIe1vMNr3ycEeTSYVmNSSx9s7DOsTKlGqG0h+o+zu5YeqYw3FpzSNBH2LYvlR7j90Qo71P
WVNXc2MWYGmXpdrkM9aIqg5yoBOyAuRQOj4bTDe6c8FOdMCf7/0WTuLz8/JTn8o1IzfKYjftLw/5
oYPKnwZpUOVogNMHzwT2Qx2rcybDfzzr8OLz7CH6TaD20R+GioYCLO0SGVvfhtP+dzurMJldYFPe
RHq0+f4vvNwk/7sjW/tg+Vx2LcPvc3Zo32xz6R85cvHGA0Czib6ndUekKlZNIBpc75DG8L41T6IN
RkK5f/OYRxQ8apEmcXbZtDhzJHGba6AoQOYmIGfny6LmNxisHVMPlp3gh6gh/rvHcJNinTccD/ju
ptML1wO/PSqDPuk8lPIz4FGG1HXcYSl+1Pz/m3qBW3w5CscG+nyeetCXgxH9KEV33F9szIOOYUEu
y4wfM0IC0IRseDVdAneRlCYEANJVWXjAHGtE7TjuqYhUTy1G+eBfvuYrgi1/iJC7pce6wQvz1ANf
D0wvJwaZkFR7pwh4zkz53yI27BLuPm4129O2sZ9YSF8dyDCujfYjiXVmrMwhApQx7oNibvdjRMie
2L9Ko2J3wlu5wCdmxFLPt9Ki5VQ0myHqM99waP6w6bp0vWec3pJy+rSUJNdf/jPmwtvPsD26KdBZ
GaeN5F9BfURbXUoRMJYxW4e7Xb6NQWYbS3B/aOXal53bwaW4W6GHLmKBcGmACAvoBC8ofsjS4miq
Uj/vqwaM4yIV57RcHzuPVnc0JGIJTGkNRfbV10GLeJdXpOaasVhy1kbOX90OT6NapYWDnU5iL1gc
jPHRrGMCckde8l3ZrxRXfS+IFvryfqs3j0MNbQ41INOOqAekQyHDYg013f4TZdbN8caTKgYCWvwF
Oit6gy8i866MzXu8fxGzM67jO0VQaXeQIBHHSdfhuvCPiX5C2yo7KOa52Uz10814Rf/lZ1dqhLUm
4Tua4ss4QgzNy5/ZomZksTQmhoYrF+LMv6p79DzUeQZGB9bIGuBCuyosV1gOfgQtotTf09EoR+Ns
qYIO3F/pKpWIgUry3oxigBhf6nmA1UWXgy1LWZgIieYRkfU3abM9BAQDYpRJG6OrhjiYTJM9ICVa
EL4tPdHvglQSVFUMuO+UdNEdlyRCLvJy82jaZ4hWgSJkFMrBK5QZLZc11rqYtmECV+xQ/4OMmZF2
A52ikMnvG3Cr4LQAvoOhnL9EfoAcJ4a1GlPkcl1+PpgEt2EhZZ2f2fMXnBdtZDOQEEz+Siu9Vhw6
aHDh1TKseLvXcDfj3t0YKbmmzEvs2sHtON4MupakhuErikv74+AZnGMkD+5B0rSJHBPg17XrI4zE
C73XQhssI212y0KaBk4av72eGZ3Tp+cKByPKjn8esMWdp3fC4eFeA6r0qM1jSLUIMR1isUqd4LLJ
c8oPcSPmIIr23I3wlNwB64IsMFpxpqXrCWNkm/mw8wFNqQaJIDFFgBWrD1lnm3dEpkOPXxuIINIk
PEJ3c3hl54tfTJ1CJcA6zUdQDvKVcBsZVxt2F+dCUsqWJNzOj01Ken6BQzHrAfiD3zG40OHPKJq+
Hk1aLFvJyWMkYi74i7pDxQYVAEdvakAIB2wkDRy4z6ymo3zs4Wa5ubeZjmucF0uuCeMITAuHuqk4
zZzTy70daR/O6DqZCbPeMb+dgZ/fEdNBbmO4m/VsHp4T8w0V5/r0SdQkwrIfN22c2AuC2rsZSq6W
Jo/01/WWYw/pD2BjFMV4gYIf1j6o/l+akM41TIgncbRLLyox57Wy70KqM2DL7sNSbOuhgQpI0CjA
+XJcGlOrUQKs7/bg0q+7Bcjb7HnKrtwbjFXqT5o/Jx0ovhIVMtAxOwB3zS9NSfD9B3atzVKrZQY3
GOsBHiQoosVefsZsK64sWHYOYPXEJ3C368GglAIEvMvBg90GQhqlSNVH68P7l6C++hPelPhRcEXB
fVuHiJAAWfQUQ1SO36OQsAjwicVxF02s6BeFr90oEfD1frdKVh4YLZk4UzzfiDNpzHptRe2fyWSH
xgqra3B7HBY3Ysnhtsz3wOQWWb6pTmUPzWixBNHmWz3fgcLvpXudKldnqubZ4OGfCjDi0t1foZRq
3YxaTI7WC7xG5u0zp8GtEfadD3AT99EVD7Hmq3qXxh/iDWFEBAsu9Dxg99vNN/eS4V324s+hnDVl
FV3yXaQP+0l/DH/pdS0QjxXjQzwS5cYwQnOzcv1PqeuIYBLQ9C7uuwnd0TAJq8YhUA68N9b1yBkr
M8QJLuAaKEcXcVOBH/j45jULt3HKanZrqu/epNOIoVSEDnwr7o42EXylTdzE28BHW+OdXsWYkbcx
Gi65yyHz4sCBSNSfEjx8NWqvGT5QRISGzyLBmXcLPGzhGopun8ca7y/JPyvKBbR5DpP6vMp/sQ8m
/wyNtOXkixNXM4ZjTfzozaFVDfg73W9v25bKaj9Dv5hatAwMPQNaVipPXjf6ZbjYMBLTu57ns3Ty
tYuxQw1Mozc1+4tE/Se/oQV1yzXbJgRoDBeEQ1rGQlQEk7v3alpcDnGOhObnMDqIObNkvRNDA2pM
gxUtd1OgfvtoqvF2BJ7Ydh+7jBP6rFvgmmxEh7I59NDhDPsbgBf6RpPac5KU0z7DE/DEiuEQ1KZl
X4rvfDGYnQ8oKWx/Z4agjb0uHvvb37BMI3igO82Emfj6jUskTIlq/wpmrFoP9yP5tLLYH+vl7zLD
HtLX1sawueJziOfQScgRiCO4IzXv+W0Ss+dg/okBEwILywUC666wZ28e5pZem4+iwAqUWruMyBvH
uyuhNsfWkjLobwJGJcFSCUe/EN788bcw0V2ZWL8IgFqDi1KoRXE7yAsBpTiFZ2sKPw72CkENhrT+
7vjlQGbYXVOJ24S775Kgv98VAm9123wAdKs7NJPHDw2DTV5sSW84QpGRCY3fc4wZOzLeiOCWPVOT
5Ej4e1d6JqEfB7K0APvirfKu4OKSPONxHJo/2wkFDimQxdsKynYJLVq4FwnO1Z5mNHP6Za7IeYMc
lp0VwQro7HowI2BDIjkQf5D4SoegKWPMku64gmkm1aZoaZFBxdVigzYz5Dnh6LlaYQNiaTczvN1A
m8vdzgneOEDGmBzAtPuGbEJ4v6Iz9ga9Afke3e67pEnKkZtV0STDljKYd3efK+9e/lEyRSUC44nG
WWivGRixM9VYxTy3o+c8vH7rBV93dNaNoecu1X3h7mBuDxCSZr3PfTjuKIatoxKB4efplx5fLDVX
+yzB5YaTqpEPZx8fbKloypkcLJzhjVL7j2nB8GGTDjfSbxS4m6GVrXt3V/S1Sk2JucpcJbUitIpe
09EDMn4xgTPgbhd9tbxcHybnSqjjzepBz/9PI5xDefOKsqF/YpEtx5bezofKAZ2DuMIY8sFy+X7x
tfTM4S5wlHF25j36BUKL0+2IYgRUEsZb0us62bT6w+27FYb5V9QA3rv/luFhsL1yEVtx9qBlqdwd
gO3diEaR0YME/rG6fvMTz0+aKdaWzNt5NpN8xAEU509hE4Dbu3cRDbpvFrNFyHct+04j3s1JaWqi
FMljg5MbMk2wmC+BHFihthdfNT/Zz3qkNoXPSkFQl7ZFnSbroJBBe7QbRI8BEfx9QVxGGe2je9fS
+GljVKaZANU8MbzJsuVsoftmqCRnVnwAAiLwP0erhk8dcQx+iWbcE5Az1zxbWyp8kPfT5laTBEsl
tEBBa0DqHD6mIUTGUcsxkPp9IjscAWzu7onww/NI0W+frxnh3rjjnukfY6hCARXQsFTunD8wug4n
ZQdD5vN1SW4ItfQJdaM34yn5ow5ymdz/b1vLvcFsvx48/+7EFk37mZzr7FC1B/ekgEmhaANUk6lZ
ZkxPjxrkmSF1DcBjDldeWvdZaHobdYb/OEL+m0ckFKHZindNWxoc8LpQBATaOxAsVH9ht7ENSONR
KaZ/LnPPGsQFM6lBiHwZrRUAOUjwU15Q3XZEPQOj/18n2xJOmX+4ocCG0thb6dzjmK/FSRsjaqaq
k+UqwfcT+Nk7pJ5ZvTrhIKinlGlSVgsYXjsoaOkGuVoAe1kfRy2zym4ZqqQkpt2adN55RbU+jCrd
GPDSGN4aPGKx3SfsscvP9ya2OV9fIgz+vdfpAHkYFz3XzoNpTjpD3bwfTW5L28hdhFwb3mgf8nZ6
Kmm25xrqhBIDzkPsZhy0DwXkOaMO3uZ7Cqz43YIYXI+tf5cVBE5RER30Bo2xrkuRGwltJAMnX7uk
ZpRAmEEhqNCQwP6YitqC1q2ZcvMEx6HIWiCHvqr80DU3ODPg1NjJ+qeTkWIkKu40XGogN+eHzYto
MTTTVzmZUZji65yZcSXlbULT+7KMscJS8eK6I0uZEBDaxkeN2OfyycXUwPZOod9R8akPePvFzR33
hECuNfazWLWrsRLRa0QOTtnFvN3B/33odaXODMzQnfeUToqKoqp7xBbYxiejoWPTETRjAw0PMUj8
QiqFLtWvnPcqQjs4wlhN1KdCLwvqijnTj4aMuANbHcGh5zHNiLXOrrO0EYXGJjISVLvjLZ6TkbBm
mPeKtzo93ZuRzYyWPkP0YGjyCznAvcDb/hkb/Xj1I9Av5FiL7sy3uQyse8b3fbgvc/PVyNn+Tb54
HH1rza+2YtQRSoIpKZfahDcbt5bQjP00kS8kFhCpDahGUFEaIX09adCcN7ybyTiuLpZ0SR5trpVc
ZsQDh0OGeZUi5V4bClhK4MpVTGC1BHyQiJD1WcVLdvJAcN33x69zgHFspSd1SdLTAO3O4Z768s97
Q/1gIjDSVu+81OQW6d6JfzzV3MLwRvp4zMBt6lw+KK4UhmO5o7RvH0kRo5DoofBHVFhyv4uPGDoj
v7+AqsWW0sJdHqZInIowv3iVOn4jHU0VdtzPm5NblfTsgMb0Xh7j5x1IdNbeAzWK0Bm7kl9iAoYw
omnHSXjcXBfxyoCw7G1f+2KR9IU47WLi23E8nqugv3oDy77lJTdzMIJbRotFMZy1zukFU6SDmARd
akN7HEKWpX6iOmf45Ay2wmgA4oL8Rk9qYv7dY2WJZYXonGqMfXRxAGdN/MPeG8R40R/1Uzd/Jtu8
GimUpAyAYk7oXym+jb1wb1aeZK5FaiV/S9H5SLu+re7bI9kMQycdSVLzX5gAMm3IM4OXtJSxm5kX
I2Ld9TCHZsZwtZA5m5/S/8WyV1TiSyf1bv1mSgHjdS5IA4Fdxll0U1RnIYNQzZ5WnfRM3UY9oOEk
yHtPPBieLDclxHOXTCAj0UQBwQdY8nNqp9KZgMyC35yWvdfIq2Ekx6j75uCKzp+HRwEeDVMT4diu
JDBPc2BJW2RjollzQjgjWQJN3E13Mut3tPxzCMa+kpL9o6jbnAwcp5xwRWQHkvR+McaTY98yO0G0
HNlo2hMVk/mzuRiL9P7+R7bbPmtvNSDhQzrrxVn6RtS3YPt0Oc4nH4mknYywmxIJ/NxSliNSg9Q+
YN0q5btBlfm7DoYJouKFJhBDWiU3uD8Xyv/n5r+4VfhWXQ6beZivZ8jkvbQDoAPt4YaOSF0OHuRL
dZ5W1u7G+5G1IYDoapnEwoEv/11oclXVriCMrSsscxlV6o9XjepsklRej11lvVvulhwhsjpoUKi5
QPxT5D5vq65I5hQEIkBB3GiDmAAjK/sPRdmYpu4Ie7Ir18p5sU37VTvIxkqMDz0idEpVsmO8gYI8
BvyAA+Ogk8+8l7ol/BvTZl3traD4Pn2XmRl+R+gzuQqmQk/wOT6GRDysgmoUebp1mM0CTLQ8zBe3
+4AfeLGvyHR+0kQYvL0RsmVA3Lm4oNB9KAjFoOKWtPH8PMfZ7A2wZZx0JL8LModxnfJgairTmH2w
OCEf3tO1ggd/EOyDIkIAAurNvgZi981Y/jjF4SMhooxDEtS1bDXKWsVKzR2S1Bx803pUg4Z35Yvf
Z/4zgNZuPH4pFn5waNLk6/cHs+8fP47oo9qC/bZTHqv61Av/WV4uV1D4MpAWmekTzvdkTz33S8/Z
7GYb5KzjN5KM+I6fYi8mo+hUqXokt2/cf+fabPhQa5pbriW6dLxjBlMhf7OfysnhQqaTG7GALT06
CBWxn+6rMQXl7UY1+3OOVkgAUCKWtP//SY+a5bQ2+s7qUKXXpWyq96YuJQQ43kqb5uQtDRwmq2NV
wqOxr/e7qIu3lm6zCSag9QzCMaB3xmU9uLV3o4ny7JdiqVTcf5Q8ODMtb9CEXOJNnnFXFVHEBdQz
71fp3OyRvmEE2i+yVWTBvII9ti5uh4sCtmHPkxVV3Z9GJxi5f6zZbEDQ1imOk+9BmMcsHo0CY0SL
zZwoVYOfTcq+JZFR5kInIk9Vqs1FzudeRXQURXUkv5jLN4rzyE/jOZF7dgCfGyc/nB+5gpHfxWUI
ll7NEDxMVXrEtH0gQjyxUfW8l7jW0ex9MQL4QhKaAntCY4C1bnooNhItlB14kmiR4NjTt0KeZaQT
6eG1zJsw8oZYiWO+YncgipnI8eKbzu3So+fuzangXJ8pJQaQc72Sctm/0xTlOGj/1KwADoj4OBJA
c0w9ap/12rOmt0RU94GfKMJbU3ftL4eWGW6hc3BRu/MHmYuL96nsqJ2pf+7laedhH0nTU55nwg+k
8a3E/zOLEOIUeYVsF4dZUAkeLBjpZC7PKtpZTkGTylWs81JzDCgiH7ei1w49a+GDN7fIJ+SHAruU
SBgPSIlXmzihWF23p6DV5rz2F/d40PCjDJi15fXXa6/o4wTMssj4IkOqGv/D+Jizd8IXIrB08jpo
B0GRMWupT0Ac89AYSJ4w67j+Y0pTxuHEmwm3wPx1ITfkCfj+ow3JZ+KoP7lkAuaUvZo5OWNX+xW1
aujZ9b4gnhZnSxKXm1R5a12rJe2G0bFWNd4Elz8vraxTf07CC5+FDsdQK+2Aom9z34D2c9Bv4Wp7
vxUjIePvpJ+wvpWwLtpNj9EkpZ2lfby3TlOJ0ylM6qtiwbFH5qoaYJxOz81nTGPYZnf6WUbyK6lT
UEeSF7DPawpbDlmJZo2tT9e+Fyt46QJSSOchgdfgjrWt6a/Ml/qSn1lsIezX+jdE/eGKkNyKqygS
Xk2ilaQUgdBnNiiuBsm7u4j3wmE8Yhhj9alaAI3rOYMQH9/6xnWj4Pj9rgEyHfOqkA9C2c05RZdD
6mF5moYrDUHmbNCAtWUInx4pWEBwNFUW3pWsY08tMU1WTwrKi7l52xAMDcwAiSHadI+92PikM5/V
yJ4x8x8KW4RESaGe5mtASY8IYkfI+MBUsngzC1iNop7Kk1CbdXOUglgkrj2rEaRtQYKB8nHM6Dxh
gt2xIKngXnspdliKTVhIxywGCE9tTKbNY1i2JDOU+K3zBjw2OR1lyphjZ82TD9MqU0AzGzWxmrZc
/hzU/eYCqPBheNdM3Kc17lgJiS6EF2/skiKSYbpwPSytcm+DVN0jiA18+KCB9sLUecVbFJ+28ceO
TYQiR9NrKwusRqPJEzK+n87+DhC0hSouX0biWKoWH0KwIt+WluiSIwnB1zb3bD17+yUKvHT1C/yK
kvZNgeX7Vk3zEBqGmF+i81Q3xN6eh/TvG9r/Ud1knymfK4topSRnuVrDqAQC//WCRT8AphTY6SiQ
YS7MSiwopZPJ8BNhOkQMFUGhqILxWvGdnjVsqJ7Sa8nGZagRFEY1jEyehYaTk7r5dI4pWOmfOS94
b63mKrY3SCNArUszv4mHWeY1roLRonjiLCp5m9lv0qonCxZhMHSTXAfM/gMGOwxnx4Igkpb5lTi/
6bdqMrM2ZBVUOEaNl6irBXKhK49qn0VDuPE6WOfaVof9Y13xZBw6fyBiQAB8Smo0/js4mB5R5sLk
ESQPtLr4+XUxLdtXZiBttDIQ9BQAGgtCZ8JsJRLksjpmQQe88nCbBNyBvZZqXv/ZlR6tUdhQMgn9
CvWZTspsq6oeueYXCbrg/gxomjNN0SvDMZeztc3MMUN4iSxYDJVuU81GGsMY2PUNO7Ch6vjGI8HF
Ow4On0zVo2yfZj2y8BS8ElJtxyKm43zwVRfq6+3i1RcvB6OzT5JStsocGLt7j/bNHFxKj28RH1EU
v23UuBFDZmY86X/4xWc6fuAzEtDnf9fU4VRE/Hkp8H2/+Xqpl2ido3wBPcw8V3u1Ny2mlhBXkND7
Y12YhX1wD/K+SuamvMIIcy0WzaumnlOBrH975Bwgo1F/W7FkmCQULlACKwKIbRO1JtrbkkMp/siY
LIdhGPcTAjiyOKnzGRYLi3h5HMCGTX+1CLnvetDKEGbNLSmL3KFq1WtzwLUfBo4ChMQ1BTyiVBp/
25s7iJ3UJDFwpgwvmcRA1K1WLU6gM+1WpZZfagpKKwXRlBuj3T2nk/rE41Jr4+xrh2SdpNM3QU7e
UpGjPLNlANRTf8RjyuJoAQXI7U46Ichq6RTgwN3XPS1jnlUkw6QOoiTWEvnIg6FP6NC4HQn70620
8vWE6vtHmFwnmjrMUkh3NCP5h0zUldIJqqrIHeqe86yz3woqB2fFSAo/qNORV5aEt8602Ji1nX1J
9CN64hU/MHuaxtwIAFHCoYdzZprr8rDeI1kRIhsJigcQIl1UcWKy+ZW2B9zswK5yEK8lK42Asw4X
/WSIbW6olnvbyd13x9VaaN+OIaDDhFKmz1BhTVgkwG0rDk8llrqgALduw/7KJda3oTZ3Zrk8tNqu
2OAs6kAFWUFjshIJwKsidVEN92rGC2ZmjgiEgb21PLJFh29P+7qPM7uwNgvlZd7Zv8jkhGHwGwge
WWO1Uz+6drKxQ9HSrzQZisgmBlWB3fF3urcfMrgiziPtKUvGfGs8mq5s4A9A/3kwXM6D/91M4uxx
XiQuJTEGnf2/WawEM+bXio3G/1mfArGOzULW3a4PQ1IxlTncaCMZh/wl1NDQ6K5G5IWpzJJo8fyv
02XERyoNYRSDmMf8ttzaCTxK1t0wWXlUEuzFSyiFnW1UsocohZp6x2aUTKTVmvibrVmCTbE/1ost
1WkyuOCgjw1g3XlakPFSxPFVOhLk0i2Yscbr/62kjDMgFtdI+87ipARpMoH7MtpXEcyN+DGF4ivQ
UM2MLjRaUlOpLaWxlWI2BXI1qms48mvPVaVvlt4xRZfJneV03fign9eJKh9bimf5Gy///VoBNv3X
a6hdxSTqHg4aV4OlWrZorv78aUpUT+2qX8kDMaYgA9eK5cAmw879EHtRpYt5NuY6REeOAHTjap5P
yzDhWJzY6aXOuSR46X9/+FJG7G1w2QinXgHXCsrjZHxWjA/AqNNzYs/g/e/UJrGTUTLyVFcTqMxg
eJSkrb7rNGyKs4NRoBgbesjp1GU3wcYtr8UJk1+gfbFVRmxX7L4+BPFTLu++TMerqmij5q9Ci/FV
R9soGM5C0eYgxxZ8t6FQZfY4tCAiRja9H2do/V1tkfGrPfEdAlJgvvnefEK0wxq3FxDC+ah0BNCP
SA+UNhqt1Ct9U7IOGtSGU70daHejxGFbElbAXEFSBvfSgz7w681xXfXSdQfjokSvtNKs4aY/Plua
LsblSovu1AFEOpTwXQELQ1x0uUv+GBWv9bag/w7wuGkrK64uxir9N2K81mklxCfx95CG4+J6GFgM
93Zl/I0BE5xwSs+LlaQoTAvs0GrGT6kwSIi99n5YiF1O8rW27YgIC8YTVdKIuy6ndfoAztfFXOBK
i0nFBJjjsB6bN/f5ZJ+k7e9uZ6OnzlsqGw+UH46HRkuDDPfY0vhA6U2SgzM7uTrmksxy9AQUFt1d
mXTTVEBQ6GoVFGfwoqwxZdtO1aXih54sakzm2ypgLVJrSW2gYyXTTmMxSdXeIExf/uBAae5stF2+
OY+qhtJ/gHT/sxfBmnan3C+qCDd7iauCLahtsGYVk3SeuTgHXQclBWeDV4hZe3tKWkhn7F6+Rnw8
qt2XlazDiqXg9BpWFPdlcHaxfoB3qUFe96JGtF5wHJCdphAIQ6Cvgm7AV1CMv9XbwbBYSW05FXqr
efVg6ALMi4+k0QlbFpAFgLDAwMv5kiVU9unKBOfR6nTl0K/YtgLrUnXAG8TkXwoW3HXJf1WsR3oS
rhkkhwbX1Zb6Zg+dNhvalJgBPeRHzYlWxUdEI//SxfNbTwOMTyNHFmf/PLRH94it9YQCOOayVzRt
gV7+1gkpIn+hIx6nAH7pU2Q/H0L42Up3fKke6Ug9rh7t1TuyvQbU4dd7VzqWB0Wehv7MirxhsoOd
shGxDH0YffueKtinGSmIXRy1Hzz1wqfulDRKYxJPhNGzzMIvaDGIJTXNCJs20hBJdc4RC1ClbY1T
8NIFolcoVPe+ysoOKw64smdpUbqCK1lXAWpbrMh5tGFn4JfRaEMdzGDvwirAjze9Nfl3ePXx70d9
k7dUWuzBoGf8k/mpabudE71lCBxBoeDmPS482FbRPtJTQbPFEI3uLAoX/ZEqRlxHyT9YnKpw5cUK
EdtUh5dDcB3dfBMxH0QKVN/JHQQ+zUw6VmP/N4ztYNogkTrDj79wwhswceBvl2NVnaeWUX1X/0Ke
gP828NC2AYUvQX9AwvhqnBiOygDAeOKOaYM6IDwrab460tFsaPIaf51YOfEVzsEr08MNgn6qvuQo
/MlEQUhg30ll4KrNwvKusVY+dTdU4NXVD2X8WWNloxRCgPxW0trsnzOqC903xcQq8xGAlgWlPcLH
UcpwfENrFtcLxXLwOfNBPO3jbkTROruO5VfbLSwjqMo2v0xq/oBaXmOhQe3vIiAVgbB0FbcPfXrc
u/3KdB70vBjbLigBMYfmpGtitIWwm8Dp3wTm5l4RjZO3sJV/OVYF77/94qzLi5exraT0W0fsfGhM
dyOKS+coTe4FoiLME4x2ZP231dobYAZ69bwab6fLCNMhUnjNLrtJnA7dblht72MDORHnNnzJxQnS
X73z3cygp46dOrU8Hdx+cbIUpcHnfITMl/9RLrszk98ndefVHoRCHDH0kgAQqUZhBhD41bweHLeB
rr/MsxrdT9U/YEqR6q5RDGa1eWj+tEQwnRJMPoq3p83atduXbqPd0umKRVmM6swv1HZ9NM2jcCZa
d2s2rqSGlsi0CpHIdg4VVGTEOAxqNRcmAVJ0hcfBDQrzJVFxUfpeCiHUT1EkLBVWzbDUgZ/A4dkE
vU8LdwoAALDEr+kLZqrtht/ghSuYcxFDBH7kN/SZIVZk2Q5ThUS4EiSI1nHgPoL9Q/SUxWhkqMkA
ED+0+EFxIfRjxE+LoixDpDp/bp0SedBGPz9lKdKhEC5YeeoHfLfJPoRUp27DKHBwPVazBDkwrIFf
TDvGlhM7JZNWxCYodEMuGDEBJ+Mx7DYTpmJ8L4kFqMKlNvi0fmbEzNHftDvdeoPL1k/CbI8lQX2j
LLrw+MU8ZHqgNYOd+jJOXrYSytSXSPyiGVBQbsmeYQlAGaSD46+m45lAwhL1Lc0XUR7zfJSlucID
9RfBUHMaLn5wrcPqX9Kf9qgrQH6c29XTlhQmniRWioR7Px0i8993HF0MoFW1X2n8GkWRrHuZ3AWH
wc+oJ3q6M/kNU6yrsPOaYaU+u9/p7TYz/Pt8FwbURA9ZVuI888UNQ1MmrCImlrFSen9yZCJSXvEj
mUof5WTEK+tNo15FBhqi0Rtf8BfqTCNCyg+m7jGPq3i8r+qp3GxV8T660D8GOx4avwM6ltrQOkYT
hPYOLItM4v5CLOy5LtKW45VvdR3CSPgPDZPJPYUS/PhXjxjYJGIqaPqW+gLYps+mOHWZ1EiZBtuQ
3uGe+ihOjgXG7KqDjWMOGdNvQg4Sv8GmXXbNGnAdUPJdkmh/FLCLdr09K4L8Q7LzTvTWyhgfUo13
e5qfTxyNB6PzvWoh0VPoVNYir+3kHRKQWJiyuN2Cyyl84L/oSb5Z31Npaf/qe2YS4aQBnxBZH+k+
rE5nEUzi61oIAQSEfMBrHvB36me9IGgt7fTOtAN9PpbfPyXsSwNjoHTBILLgdkOEFieFwweVrWhk
pw+4HWzZWM0e6rKKkWRhoEOEDwvmnwbuHJ0J8sBocJDHxBOE8jvYXuIeejx33SkiNptOFTRW6owt
rZhLzfEsRdj9gU77dEMDkhE0r1UHjLSe4M3k1iii3Htu2VKKUHAnHJRipEDWGm7BncmvXVhSnCGR
nyrFy15wPJSYJud1pqgZugXp4S5oasLxaLqR4DvgRdGsF4qT4d/+V2mQvur18pmrT3i6QG18gLp3
krUAYO7kka2NDEtqbM8/avu4z7QXh7Iaqrk0excW5WIbIEq05L0P1wZUK7OZwdaefnFrvL+a94gW
+8pDOwP5Zo+gM5y2X1oAOG84mYk2/DZl7cYxSh7dGi9ZJo5UBbYGD5B2dH5seZU54SSjES5x7oP2
xt8tSE/WdQey2mUVJE6+wVlvkw8KTFpyXtL5+jvPnPIBovOerRAtqHcZkgPVmquo3AFc33/VWzUv
K+H7SlLpDM77jyH7xZqsB2Ht/HfjsE9yJlV56KjlZPT0m00TTs0xD8vQnhJMv42OgEa2roO3M3vM
svsuLEcfejqsKG8HKK7KdKS17R6CSz/jCe+8aMPbzh5wZ5BEqdvz4Mq+NqS3QmlBuwSTCSmJ8yvv
+GI2cb/DqtUyFevDU2U0cw8cxqjECGDDtLKuA/s+ydmaY+s0YIij/f6J29MyHt0LfxemV3s9sFoC
O46FhzsT/9rFbE+skIoa4WdmAogkSbGtFvmQayRNmFBpkaElCWXGA4JrZ+A/ORTXrDiW3cGP4wpH
btekUNL0jdNGA2S0ReKF14emH2fpVsleA8iy52mia8MUWlBoJZwl3XbR7llypuADSViIXfn+ji0s
GRSnYmRNCqvpFx9jmg5OawUy6SZMJ2URg3j8j4Zob4RsXyxCYuCdWcFcKGN87vzToHJvM5gVZpet
LDIW/1lW6x5GonQ/k/Fk8izcxVVzqCz87rsoZFJrhU23wQx6VMDbBQ1NGN5iP99/bIs7MgBsL4YN
XkfoEfh36Dn8l6gQcPEyvASSYKLwQBwC2do9mtlVHbD7rOa6/qa6v/ybVhpx8TRbeeS3BCrnTk4n
oBHciAHHHSBK21dgiHZfncGtsDorBh4bXzbhDpQZ0cG/+PNLje/O0spkxUOppbxq2e1aaNBjoole
Ky9lRsv7SnVvuHrN5lD7zvJh9UMXHljE7bydzxx0FuH7CjvCahqUFa5qMWgqXoqK4JVN6sMc7lIs
6NM5GWcnLmJAWGrJObsjNShLyY2N9oXBqi5qeyCyBvdkWsmVThVjxufNZOWbE/hyb1HcSBMpzLTu
pImnjfVA0F7UABE9WvdhaSzzBOru+MtwMsx2HTsQW82vjpapCkKVHxYlx/xGGFhKHur0AFOTPyYz
v8bR4fHdi3ZGEn5J3JACOkw9dwQgldJJ4gPkltAITW9R6F5gYqYaLtePIFxcZ7pVNkpS6i2vUT7R
E8I0Wezu+CFVWpeU4K1WpcoAlljH5odnQFFQNAUXYbZDF5/GLpqZbep7BX0efC9TaB9+76gvVDE5
k1Dy5qvjaLcRH5mALTPK2to0/WcaDTeteRY2J5ZQSuJSCuDh2yeVczJPnUBZQwpRcAu/mEoSDEeN
OR0z3RlOWtgvnM6CbpW3LlOWXV/TYJZ50D0rWPCg3ytbQzrINvrQd/gUxtAKaeLclS68VJxMsqLG
diDJ6HZtKz0Z5arG4IEQy+0c/Taj4/QnUBDpqCuhlsXCV90/+0GntdebPPViYH/RIzO0OjVm9+IW
ybedSk3njgVqW9sV9rTxVuU182xfT8SAAOgU2S9rbvl+UjV5RaUO/3TdSJlaVPcLbBI5kLEm3FEw
RJbUThZCU2Lqu4rGQf1qcB3X7kgnKxA5hEcEOnyvZW3Mr+5AHom3bbMBBe1qo9fcqG1A8B41y+hN
zAdXQNle70XCtBzGF7QDhGmNHw58tvm/LBud/UKVfMm5eTYCeXdoB7+/X+Sfj2shpYbjMYaDqTx5
NpvUJCa8jbgECPUhNnOYmLhVy70q5duFXEFuvm/HD3muok6i3pVMWaDuYt8u7J2dv6jG9Huun+eq
3HICvyG8U1MpL0YeDp50DEQP8a50yx3uHVidaMVLfQG4Ccr7sTFDX4ui2AmVCyTpX+16f1IjSGl9
WiiT17+oQs7qq0oxK0XHdOZrPDDIVcmzm5LzncNaFTvTwbMp8H0fnqmEBo9j7rgGOPlzv0iDdCt/
FQTM2PzJJc2OfxvSCwM8DCqkWRU3TT4NO+aCtF+FS8U9tFuOfLsZSIuoAF4SsldgNLrEOtUQaEc2
sD9DSQWK6xmnwOwR6GIXjpHQ535FQitbRdVSRGfX0T5Vfs2oRs6AjBqLFSndwvFc9JsGOpzv0mwP
K4yaZ89GzkRustNhfF7UUD9hkanxAbkz9Td+V5RGKTVcBsal4fMfT0UYh93HixUcymxx7DHDxI9A
XCR80VxLdqk0BCiALqH5mj8S4eRYvN0nsaPtWGtTa79VYRTan69vwapg3tVIdBw6OnpnkVwXfwIW
pvM7Lm44vJVrlK7AgUFiQoNX46U8VRlBIQ6jfhxiuRKIYk4UUKWPed7rKoJMLNLakq+NPdrG1PXC
3WpXTd0+Fau7LWHjycayRQs+zYdlv1mvQCZXh9d2HXd/BifD0OW76Z9upUEktD55L2LZjHUGjgOc
uOZPHKwUS+4rVqa87JImSpl1sPRa2sxzzaJwqXVyTzC4vAqndzTbieINFVmYanwAGx//x7YSaWDb
t3S1W0O4oSc6zT7dhIpHB4Cb+6s9VeJwnl4MKvJxx1qtB/Yt66CxI4k2Uz1dXBBy3L+6JhyTrxoi
R1K9XuRy0cur/RfyEAmMnTjiP/9PGvAMbXbHVHHHo6gd6vZI04OsPhP9oaFbunHJdXQv+PHZYZJZ
m2DJ3E0JROTbc4TCkAr5eQUeq/vWxG8m175yCEoNE8wuGyk/1j2Bzp67kUeV2OMFr095FsO5jO4p
0KzX3M9yD1H5mNpiALOTtVt+J9nn3gKeIyRq+FGrb26pbHjnd8VX+RqZXS/MdWITOjHxMwDLGXAJ
Jv5N7zgkd93xy2pgKuGVNrNc++JTRk74HdWjbOIXWfJT63oz24qIOFea//3e9Vdg080F2X+2j7Hx
uENLVZiNiF0uEJZEIUo7ifmF8tcmMzlPg9PTvOMe4LRTDz06BRh9Y5DGrd9XlNhaKghhdLgLf1Tp
bpqt3OLhE90tPIyOzpYBhxOX6I6nrLsh5qhK0gPu0xZwX3SFsddLM7olS44XYsyXVIBnNoSTlp4h
RyRyOHHLESq2gDHehbEbo5Twjp2Btekgq5ySFhXITdG/e12rX5p++UOvY9apWqDrSkCbwpNQIFk9
kdThUDrySu4AC0wTzxhgPd14MyVgpRwsrjsubhOl5hvBvWNvW7ABlgEjdN2/DeX2Oumsp7X+858r
Z7Fx+OrdF4Zla8sZKRq7zvBRerVbyNIH047ytA5qb/9gmL3YlbKdNggKP0sgW35hH3qrw8XfDo/e
xOpElkvRbDf5Feuuzqw9V7AyxQ4yU8Ht7obeN5UbH6Ph2NKj4b0cf3S9/vs6l84hlFpkUizun37T
4c9EtxDTAqNrLI11TiyavRKcCRGHKJx8HsVxbTYPplAmXKJG/Q4RYJaw56799wMoLGipUXzpzXFM
MM4MGolUrMX5kmrcqV/6copd7xagdJc/BqVDHr4OuJ7YvAB450sxioTeVqWZq99+/TWHKjXceAlG
M2csYtL7KAQ8a7HrbVFqXdgnvoNduNANSufYRYAxy4zNM20QQFi0gNtNehhIjcvex51dpKQhhC4e
v2+Ga7SXGhuucMEIK1zkCmDMGO1N0x8QtjFCtkwCiVMNGveQwjt4uR55p0/QvWm98tnwa1hVF69F
eG9eC7VIGcbEWpRwaLWK+faOpHeutfQSKmVugjMBPGBu4QGIJvFEx7kud1uwjm8XLYmdkiWfOPVa
oVZM3Cgp1p8a3OgGexRXyWodLVQ9oprjbdYIL7ugjly4Gk3cDp3LSSL4CPF5kTw3o7h9APzJM5vC
kbSQclQjapv/7Efz0rOqNCCYLo+7dchVh2dLXnbbuwhKElCSQMHmej9mTjCKjMNeSvPlKj5755Sc
Hb3Jw3hL2MDBlV/qEN5pVJzxx7g1jG1kMR/zP6cxYCx53ocmeTz+RwHg8JpbmW41Yvqhdbk2UkNi
5G2u8Zt4B/EZDoooJTWbHHRK09uSqMLw0buwTU0sJT1qCKaOCR1o1kJgej3rxPQRd/LhLJTYooZS
OL2fo2Tstm1bFjZArGa/7LiSBwMdqTJjYhx2nWqqey4MZSdp5UEdLgB+ug5uFyT5Wd27SaOFjE9S
IJqAMnMnOCBk1Uq26pKUlry/gqsHmLoP4jE2BwLzR/lnjAQlCcLwW0kosHb3NfJiAqCXdk7yiAnX
31umEQ24QE5ju++v8tz56P87JgCIQ4zCM99NAenY2z121vj6FtSZzBUT+0p9s28ExDE6wESouuWx
oHbZ1re1ztNSdZ2CXV7ASSX23p73j4XHEpB4cNw00/tN+h/LHod6GZ3wSRDwpE7SKLnJzoTqj/Hu
EI2x4T6ERl1Hxe+Zj76YUK7Yf788S1cYTMGTEf0cwD/yLpJhZfU+YyCCi/s+yQXdVX/pGiW5f301
SyYx6Dh4Po5G5lX+Z0oYB0Apmroct2B6BEbl4Hp2e5FrcZr2ueQy/Fe/cnh0p5KETr0IKMmD2o3N
mh7wBi7YoaHpjbCp8LnSxmp8X15cPn6uQ4BBTMOAslDx/JPlBXdlDrGropn2o+yD6FEiofQfX6/7
CQ+fdpHlAWbXY6WPsCti6IV2XbuLWUK9oD17MoLguagY/pq/MOe8ewI4MlWVxw7wMaf1gQAHYpaz
zQ7mb9rbtT+O9Vgs7ShzfNreodKAXPTHpDoD8YECzP1115sCnjkJyuR9aXczsIvzUzqDPmmcpCd6
nUBWbEcFaAy09Ti6dMuANDfU6HlYBvC8nviWaoq1kh+Dtln7w/0Mw9lTd6T/3arY7Ix6hjJpoAzr
xJ6AkciwI3iyXTEto+cpf23piRGeaObfav7gO82yli31FLkNEiGlXsw77RM3jpPN66KfNJO4mY5z
A1hlq2kEx7jyw9hTKWx+7D79C9qnKRJ08QCjJGWeof6MyIJb2xUg422ZOfy/Yur3//sOeFfOEYIa
FYI/hK88NRxjxX8mEE6/jWdozeL8sakXmMqbo1lmkX3RW0RJEA1wDokvGenxPvxiUreiWMgjGLKb
zLLnMwS8wyluofg8iTvsuZq8AnoR55Ni/m0HzfYkl1f1kF5o8jPz3uhMS2EDx/sDxerKYRrDAuBL
zzhJOkldYSVeUZX6di+C/RnDkyR8iwFcVmqOpwNg9fChXb7TdsSzcDDwkqgmgVPfs8t6QIV16dw3
NaT9iUBuP68QseOOpXu7zN5CJjS1s/I/gv4lZEJ9I/Uo6ex3Bu2dP0JGn4mQBb/i3Gddf0i1yyu8
FOYAsVZoa3ZewfPyIGqBLfhIairh8zwnskcfoT4iDnKqDG3Ir8lzoUwxZppg6y1fAontKcFVoDgO
XM1VBh7ISdU9aevN3PKYqmMeOsOiA2k3pdzGkxZ5Z5usBm6NXBwISWGTocQFXWBjixPybTaUwlQ8
ozZL85OHAWVFWL8p3AYs47KIUObsprB+CQTL1U7Abv+DIem22UUxpsRslaEp8eMGzQnKivcOZIbm
9RjObCmfQB2IuoOVNs3d5ZIAxZ9asUqDLmKpxznBHro3waHqJh5ImI3vt35WkYoAmgBTlgcYbMk6
tq6/QbtqAeSOWuozL+orhOXuBOjq/3MSewO6gXo8BOGY9HYo1b1HvERA1aywyxKi7CqM5i2VbA32
x3hnETP8lAJhz/kLcwB8iqpYcM3GRdMB2Q9PxMm7Nu4A9ueG4ZNgAvGVrso6ercgVkWumHaxwauP
LdkYJv2apv6zduDwgw/ZVmsBTLg26T/gnTzCB+g0ubgMQfpo/Dh7P7+9lp/a+fUJNUFi94c+3cvx
usTv+O85vobdq/7G+xbGGGeyS/CqjuG1p+1Oys+bgrHD3Qm0MgsqyYDie+D2CxVAyBEnbHUcuK5y
XYSK219QV2aIIG6J84oAhRT6g7iYeCRv13eJpWqv02/lRsT7xPVEFIipSooXL0YDtwsqgP8OsXHG
Eex3YGwsiuIYcXYRkD9sJ/wXHzAkC3d9Fd1TPE82KCVbz2LTt/7vZFXf/nqatIxiR6MtQMKXCa72
WW4I7dJSO5w6vCrdsvGvDibNv1I2SEHuVj0wdxRwrVYp0XRXF/80IIIOJPnNVuEmdeba3cY9A25R
cpdkXLYrTXl1GlU2fDaWIhqD3lR/XFtNfyRl2EQScp/Cf3tn+OW1SNWaP9VHin9EL6IOtKB/N6OX
GIXEFxLYaHX8qnDBmTrAYNa3A6jtELeU2SqWpN1ZbI5TVxVBBpM793af4Ml2GDka1qnNsNeX+ujZ
F85gp6uRURaUxtFH6srDo7Tn9+gVsCjJ8fxMM95xRpztm3wMpWtl39nWb36gAg2GbLx9t5GSdmeS
t9GpGOqa0WdJll/Wu3bevePdea1eQueJD6f+8h8E7RFzU4GKDNwCN2EFqC0gFPO10si+z0GO+K9W
V/rAWZCRAcMFoElTs1praAjaojuqqXwYenrDSKXAwvXMsTSrfWvjFeo1FzBpMLXOjkDyO41/06jy
hWm4lHRSn1kCCKvzHpcC57b9385/SSjSUiswbnyp0vT0GtgZugEq4SaUAndeMNj6ZtXGv3APh/ZN
iFFrILWbIBOiG7Zwb6SO/aPcgYY4OFe1215rNQ2TSwOVTGKX2ZLeemCghaUYcEGBPHE9PbtQUU7H
jxF3+crC2yApownVlu57pFff87wJLUEdMm4X3MxJFWG8OzyXYte+PWB0Q9BaOt+qruH/PyPxeYle
A5Ye6Ko7o17svsekH2o+dJi6HYSWuw3e93wOcB5+Thn9l4vA0qeeT+giBENj/u7cNAJMEB6w1E2V
P0hO3oulpNgAfbJuB689XKLIJSkqoNZB3e0dcVaY8zuVtBQvu7ZdtMdwVweBWURm1nZjY/p15ijA
mUU0HrB9NM2KVJJfMmxGD478xlk6VfUlFzVZVrSql7OG8BD9vzeeFmZzMSSulUV5+uhYnnDurGUi
CeNOeO2wl8ztY5V7QKME2XluZcpw9Wp5MLjxcLNia/i7eAQ10fF7qXXU3qaN1iN58u30iVMAts8h
JCga8llhDRM/PCs7ZAKQODeBx5oyYpQx8jIEdtIsaBC6kbdqWPWbT72tHuKY/ohYa0MBK8RMLFQa
Za2mJRc917BtJnhyM7FRe1U8zqsX3sxy2hD/lH3cBls2iinLrQVNaWKhaQg3a/Mas2YqmTJxr/Md
co3JTHDmGrurPOmOIBNrZ50uClkNik8bY0owlOSTaPTedUZo77kmidjN+hFtuv6tvwVsVGL0kozb
jRgkWL9fu6QR+0Q3TL+wicJorcw6RC53jixu0pibtlqI7CkbTQsZKoDiwNWQpexJkxG4IsY3pW4l
ke9t10tRTdkkQGT2ILkDzi9UBU20lBsESPdDdRQ27gj5MYiSjQFoHRTXYwTeeaxHNAOqYdWjsrLH
SKIzn6ffqf23widm9KdSuteGhWywVxmuJ9rikIlTXdYs8Q3Pt82RkhCbILWlM/uCVhG3NGuLELJy
2+aYiDVXHRJfI9igJci/I+owCUzFzhM+uT6XDvcGTfq/vMY7y3OZ0xGwjwonumAiy6+3j3UI19Cv
yNnJpRGq839b9zAnO+GGQN3+h3qdDn7qZIhY1h8XWmL5kPOEeT20IvhU2rl/rekwh7lkL2nHxG9G
2FPq9cIUfAJ2EEih0xO7OMXQVwcuGYKqPh6ZrgJTDge94NKYL5SIcJQj4pHmjlsCO3IiDoZ0Ow4q
JZrUHzGQY9i0DyBZTcMAoB8xjLArIzNARKQEtWNAa4OoY/AvoHdVo2RYVhTVisagWnPfADRSIVNz
1pOau6pvNy7CiqiVilefB8q2YKNknoZB+m7GVPA++cocg3iYmojjwxcCbjZRUEeaGerSlgasequN
RAgRxZ4g2rgOi8BpSQEZYoPejrz+/xYO4zJbOlCyhscpvAUvJWWMrNvDu6pYP7Q2nJBri4sOYOnU
GIGeZgywvRdfCGXXoQqdDQPcWNtIt9c7LMok2Hc/pGvWhIpuLx69NsuVDSafkOyTQcDL8Cu7a/Os
JhQfuU/W4d+0oR3yjD5K6EmS0cpk/KSG8mDB27r6TI9915PfNCJaDguhTe+5BnCp814nfx6IcbpJ
BYWcnUl+NS13nJaqmhj37Uc1nMht+hOIo0mm9nE7QOpYXj+dmPSPUkLvunCrXx0IjqTYNkEgXPsw
GagHcRyvdIdtFLb8RcDqwRqrF0H+NEGlfpedQ44hhIDndgaA7kp+hOPYrZGY0VAuQAW47Ti4FoEB
PnhGqFpk7C0Nr6IfO/3OH7IEzEmii5vAUsWh+6stzetw4J80cAUMnJHOyDKHMLEMYfbc9Hkqsu1H
dveJbwAaAjik5QclLNq7lQ76WxJmXBRP+l1fv7WKCpBAu8Gz3+WmpieYrY14U1jmGW5SZ+k5kJLl
UtY7fepofEAjm1eEkgwGHCQwSZ99/aglLJMHQTLCl/FOi+LwEQpQ3bsX+f0Qof+TAU+zdHB6qmid
9Dbp3dmne/eV9g8batmFLwBFRH3/rsqP2+1x4lJz6cKraNCONuo8LbORfXL0D9GHkMPd0UME80r1
pi+rpT2tGpWmvCwKOLU9j73K6VGRoOVcnWvvhPdKrt2eg+MjsnFAWCITs7OFy2zVvk++poGWDLWy
FRY9R4r2iFJU1WXqQkF33HTZm+3Z4/5eL34uZcKpddS2nQedQ93DFTWEdCxTh0XwWmbY9EXnoCMl
xeaUQbvgcirUiZ36nYX0HeSeMam5SMcfW9Ss6G+ul7Bob604uXLh/9AjbS3a6KE5pyrqo3Ix+lwH
vXpy4HhIVr1M7gVzHxumfTZV1u1iwNLp8xLuDPF/Sqgw6IyJliQZUSl2US7oQnE2kULhsI2dW1Z2
cFxTpL8jNCzDzPm0mNQo4p3ytQlOFrn4tPMdcQ1F9OvRkOSn/+peUPKYpZ0+FJtnxKpJM0W14cGN
1jV30aeVXIx2KJ5uBspgLpkWQsBOmFogZLD+h/HGLTDqzajjjeG1J16dEUO4qxeC1SqZ0S7gLTaB
guYDWpVVEfN5Pv+yW9vsdJbfuXj/1fRQfIvKkWiV/4jLFFJPgiWeymKHFGttHyKOIwPpHvpIP0UW
PJMBVB/CNzOytYZXFk9ctayobwbHkSdWp6vInCc6iWZgQsNTfIjd7bpn0HzMiFjL9MvEYBp0prw/
7FpMAh01SJQDU6WpAXlZptoxj9oRkg0trKJfDdrsCTnGl2Cv0HhLJQOD9Ozhypx2roNGckbzvGa1
QKqXZJli3nDV4nVKkp+jLbHDlQTqT5iHaI/1Hg00l4d4sG8YABKa0ZvUyP7TB1J1Fmu2WikK0oT9
rPkDqeFYY8PpI/QZZowtiY8U/1AZsMwavm/Vhws70DmgFLW9zIytlFByrCdA+EjshH2H7mW07QMm
0yu3PrV3FQ1Vsau0n6rzSBYuDLSW1OKLejlmRQRha70C64Dcmc+nuR4MChp2i7+kHzLqqU5wpjLP
E1lHVln6DbISyAtiKfWxCsrgeMy737U6kNMsRBI7LY9bw5Nh+DJOSZdXyiIOhbfJEt/fdaKyMt4U
4NeKw0hJ9wvRQyzBO9oq/xD+5aiSX22Yw3+MVQ0K2+Lp7Q4nqpL02YXF5F4WDTmC/KQ4mdYa17Rj
H566tn8aLk2BF3AuatChCclUVC+kWiqYTx5loaTCxxO49x/GZGlwhUf98fNOL9Py79VMBhdQ5UZm
E/t6mMsUYBf1jyQ3idGWxXyHsmBjMaHqN8HYVzktdnJi/DMFa8Yma0OdbcaDekQGkwQessi+Nelc
5r1EVbwbCD0VopeiaxM8d8+WQndY132bjNOd8gFiUG/z03F5C3E18rVmO43TkE/1/nNmB/6JAjVE
uHczz8JpSF5inUNBC1mqf+K29/QsFLK65cNL6VrhSZgm+67gU0BnTVJXl9061svtknBa5ToanrQ0
XzDq3vaoUYsy+efSMs/+o53oyKQYou0twikx7WR6BlrnOD1d1rDJbDBzlzmlK0GD8XZbxsNCbI5H
oYZZ7D2arAt7gBG/zxJOsdt+DRG21EPFMxBwdNdYla64CStYBBIRiagFnWm6lut7l2mroQGAvZ4R
B2d2J061c+O52HYKlpjfnHetJeA1GhBF72irVaohLMdA4xKDnWV/UNXAM2w7gdTzGE98DS0GeyCG
B5DzHqR6RtWYUKZzusFszoD7adDrVer+OW8K8EXJwCoD2b84OsJHyXPWePc0nRTsBPTkqtWA+YwK
wB94RA0c62AhPZ/mieT+9UotLrsdGHOUXK1dTLjqP9KYTNtM0diMzJxBFcMqBLcdH7FvyNlfygMB
q/Ct9GLA6zv7MCuaN3p67ZNRDhkd/+wJkQ0/KLttacWll35Q6ZvuvIFhKlFmVveOYxDgnGvIdxBw
bayuwgNQroX0Np34Dx1J8cc+JinRblZ+NxwqEmMlHTh5URXAhGRJ409Oh0k6MeV5+GzU0EyW+pgb
PkMjElUJZc7F5n6CmGKzY1C7OW0ELJWyPDraswlNAH7j7W17di+PXWpy9viTeju0aQbhy8toM982
kfw0zqovX9om3ObSnlIQzftQ0IaP0qJO/Jn5vhVe80O7C9T5iTq951rtqXUH1bp9EoA2wOTt9Jj/
7dznZnEiW7AkbcIxPoQJKk8CpI3DlxGLQbaH/v6c134kuiEb6WLsvOnv0nvJUj9HkdkzWYUTPAiY
dT62Bg3Fgt2FKjFjVMU7XNDOecszZ3UXPrr6+DU4HsKT/cs6gqDL59HUO+yxBC26XEZMGtI7hdZT
h2e6noA8tb5lS7dOOKBggVjl2AJc5N518YHY6WgEQKg22FY4yWLxV7AIm92rzBwdm4FPmC34eL3c
fSO7NjbuN6PM2trl/Gr99YwoOq6VzF43wSwKN22HQJ9BQfWlomj47ddmjKOZd/sZ+igQazoT3n+Z
C1NQgkLe2UMXXjU6Xw2LDJUNmrSmKj4JZh28UXSPjb88tdPkTXuP42qUYO+kS8pY/UTMyZummNCD
OmI43LEQOcda5bdCyI5Vb3o41HUs/L8UHaYuEJLhpIOr6jv4F6+FxQ+YRAC3pvuAETkETY/Tg0Lb
qhICMTCLAUM/aSsusS48XpQ+flZfr29UkKr1GEmA5iMFCnzEuOd1u+Pm3BaW4pJnzhbfy1vm4nZ5
oFEVfp6IQOsiWUMQmem1ICOAvaQ3xOq2k+2PTCAoLQS/srTBj007TNlmYg+dYRLe4vbMji8Ak/Qw
yHOZSkeyELLywLASxwLlWqj4ooZqhvX0Aqr2G4unZfT+aerPZGDU3cBU7mTP8oRx+BXM5mSV6nmT
8CCEFhtr1hlNXFUu/ncFDbbyRmFFV3EPwJlphJAk10XubSP+x4VNssXzXwdILWWu+Z359EniMZPw
D5xAFKELK22uZtxGM1O5GcPTIVZWtOz6tCkSYQppC8pVwX56Tdpa8OmoTn//4bYrNxSTEaKuDlMx
zH0I92OpjDIti1lWR1m5QEKkU9HTYA287XprCXxDgTvaDIc0TmxLZ7sGXvahs6Cr0pBEmYBo9LTt
UwLn3pRyd/mhCOmyxnhsmmMNXOBsU6MljyCsRu+LZ44etCgenhfLjeTk7lKNGBpQCVqZaLXU7ZDh
Ux+80nS0jA+UJRGm+t6N8O/e8p9hUBSJCXg0pWpTes1J9bAK7dTsb/40hhq/p4FgwgRnw80T/bFM
QpKVqXKX3GhBRGO7gggcgh5+3izQZUhnCUYqJzoEuJQUy0EDbyxdKBNPOu1sBpQWUEUP7OQ91FZM
K8GwqYFe1uDT+4PiLXnWTZ2t5oQULbu7pSBVmq7Kk4dYqH9S7FEMxJ6mq00Vl8mqjK4SKdsFr5XY
oqehws+non1I2JZYPldHmWQsdOhju5XtycVAYz+UDMgEfiG/jX7eY+ArUT4XZK1bNEdp6joLDyKV
GdxV5RneZrk4afCR5fw9R2zxf9Tzo2obPi5lVmLNMK7dEZtm7ugPdyapXQXQ3esPWVNjesEbwdJb
6o8SQh8G/RETL4w6dhXuiluk2si3VsBv+N8qCv00VnZziCFQxpn552fT4Wf5fJXU2jUkALiOCgOH
/vEqkSxZV08BHZC0m/vJSpq2wFsIj2rvGOO40sqNrugH3PbOtbZC4nEE4lKVfB0+/ZlIC+8jmXsa
g69Z+F/sceNXiSGedYYAAl5mvDNqQ3LTRVeGKyDP4MOSjngYVLdW8mlZfhxxLTBbsHDFe4Zs6oXJ
buOnU5YCpaSQZGeaP5b2jpY/3Sm2t3VGq4Vbt9SwBzDM2GSTjC//UOV6ncWeRBzuvqZBbc8mNIDk
JYHznh3Vz4DBNttb5q54o28Wve9Fd+IwdHq75ojgT7CTXygnD2qK2BeatJ7iq0D86xtZdWh5W+WL
uKRwrMPVV0T6Fk2eZBFwFRVRGFPx3HL5T/Z94jgckIvja6AoN7P6J+iislF3gq9zw+GTfsV1sFQT
aI1u+vqNISTHANiC2FVL/JvGeonV4mFb2rPnzlK0OnIiTlgx+/zJuVv+WzR6GYOlr3UpZN0L/lsj
xSsJ0XptjP/08shpX61JQw+DiXpqljRNS5aE0Er87+UL2+KNgEnKiFnzVyfkoG53qQ0D2arxNHcv
7dki6pGl4iAFdPIJWyoXiNycMU1ZP7yap78sd1KSP2dyKARR6fvrrrqF/Hp2+jk8bNcoAD90HtqW
5oPyPBk+HDb7Fr9WSGDEyLTXZZdQZ3B1pJ4YTsoW3yU67ZgVn+dseK1KVH1IjSp9GoNz4zpkOEWE
mfM34ItmT6o51mQb9FtCYV0WaBPK6eYf8wVoujAjn7Md3dXlz6Lk1kvEQR6QJVIB3JvphNkyqcoQ
L4ExIcu9a06bWCVtEuafpfTO4j/JqsLHwZ+S16HjEpi6s0vKGneEvPAF5FrIprYZxpsdSDlNnpDd
/bX5vPlZ6qAW2nCikp/+02nCnwQTiiJqS9PT+bvVTy0s2QoP2wV7gr5bM5EvQ031O8j64iTZ9+Vl
RZcAV4HjyMQraMQ6YDsqe3s4Wy7OzYTLluWkdnHRgmAiPxnoU98mwUfJAEJnfyTUDDQmTdtYEvht
2cA6k7PhcQc1tbgGCJLdBjc9TB1KjLdYdzWkwlI6K6PpBJhcJeLs39giGDvX8v4IoeMGj+3u8MIH
8TshicTBXvefsx5UjD8zNbhhCZh4LBzSsLhMtfkfOXGW3NsBwrue5t8BqPLjtGox+qeQV10lZCKB
7092F6iQGkewm4WxxErntXDuGMD5WDE/kt7xuM1OE3g4zlo+2+4mXYWmmB0Y/Lg0t6HCYDHBWlfo
EHYB7RDtuB54gfgZhU6Mxk2i+jUg6XMKRS9AdIXWjj80O1kRd2j/sRGUOdNfyrCSresF2jqDNhke
0JXS67T7+ITbomAcktryfGDMpg37W/lRRfKheJ22QpgSc1dmEhCUoLHQfEY5v6y86rqXzwtXgJnQ
KWJxgSUkuYosSf8qpvmMUuo946sOELmQn8jsc2hPE5cwCzovueAIqIUBzoDVpm4REzfQFHR5qDSh
T7IsCIA2Koc1baAvdnkIWy/rmItHFQxuYmSAPTjyndZHcljddzDchd791DF2I/LFPWahGfKsfwbu
l9kV7hGShB/wYQDsK03X+ZX4VKsJr5+RVL+Cur5hSGROHiS8rUwrZS3ylo8YG1Y1elMM+SlYGNuc
aKCOpn0JWf46Ft50XIjpA7BjFz/a6CqdplJ208bwcv4ry7wTDoA2fhSHNwDnQqNxZfIkkF5gzB/c
6zJH9RwQh/7+S5/FaI9RBInYDhvP4uhoDE9B/C0fhRLzUWrx+L3eHalhUdvd/uZh6lJRgkO3BQbI
isJv8tmGDqZsBoWglvGQyHXPCEe44nn5rzHHd5BOebcF7LTLcmWChvAcnOsCm8S7aVrajW5QvZiG
P1ic1wP3FVAak4aB+mKx8HaapwZHjKkxWUMiLhF7GwsKPXpo8cYJn2UaRDPGvZWybZdsC56CoaUR
x7I0IkG1QVly4RPlKLAaL7lLIqGuomNiFXld+QINgGP5UGMjUQv/nPmFH4qHZmNu1m4kbRT3aCqp
n3USjrbIf+v+9vNOLmu7NAGvMTIhNq0kRCiVis4YKproRlukZ1fdSvMXoQuOv3AhVYdh69g1Qf/C
FwUr9+l+E2HKGiJbeegr96XV3C8cCRs8+7D7lkzVUQHmHUuGdBGG984IjVw6S6Jp15Iad14EHQWl
AzouYouJmzP6daECkaSmV/rFfoQB/qvwjQlCEmntzP3xa5+2Yc+NoNbIPfcr2iWJVm7rlKrD5nl7
E++IDSlVbnpNZtuzVl4nxjuDZ+ZHGONaPhy8CNzcwrqkBKOG7pulIURk/m1DonreqmVzNq9sUc5V
pvIu7Or5AAdaUCm+w4CndNfOyyw32WyTLqhUeabL7Lb8CLZJfjS7ZmvLBXWQMU2u1RT+O7iDMi9X
ZdrzZMm/oDLWX7lwXGDY50bBOzFDRR85/x/ZolgKntUAobGGhwR2UWcV9fk+D5R/KZcZ41dBgD3g
8O9q56vuK60rldI9+IHxofEg5LAtQ+Rvz+q3EYqRgkiIxWjNQKNO13Y7t9Z2mQvWdnSlYyJ4ZKDY
vXIl/cJZTP3dqLdJYckqkzza+9QFPW4+H4WnTv8OiLLynP8UOSwr0MBsT9o0Yfw++IZgokMlBNxm
yCdy7YcAtWESrsrkmOPpBx7htgNLNIK+soHl20HZa/1QwLjteIJrvGVnRfWCuLuE8zQ7VUVTSoen
tnn0MrCqSTQ1xh6VcVHGR1yU/rU0Y9rVD9G2Gh16ARL0aosz28cmSmkRaruEajGPQwxzz/N0jvw+
m9X3Q8vgOa1Qj/eQAFnhknatKjXaH6YkDI28uEq6CeYMoJrEJQ/nbHyH6J0RlgfG9Iji+Nl+pfLx
AhoGCPJmx2F4QHGKojiVGqS/z+RrdIhX/O+/DPtylQWSlp2lsvRyTCQWBVt32grGWBnUswd6VO/3
X9c9nOUf8pKKgzpZ40cCD2cv1X4MD3H/EMqYbZK/vpWnsX8LLsRUmbSp563M46liKAieHUo6MdMy
WdOIrrU+PfoAkBFtStqikFR02euMZiN8rQlcByCB+I6btFfJnTgNj7k3a9ImbhHS9Y4Y/Y9kAWc2
CVRBhGYazoAuvtpGw2aoXDt/+0cKELrdpP5QjWmgYn9rpwGYpEod7mD2H6dsE06I77f/Q06tBp3R
R6mvMTMOIOw0Ynt1gtITfJE/4Nk+zv8ozQIWZ/d7lU0+mVhnmLZlxqENPFa4c2gGYD6zrPHEFUho
j8ctGHE5yU5AJLYpxkiUiBpwZ2nVLat/WX1dCpGq3lCRoyQ4Pd8uWUwRzWZvwMmptul54EyuAIdj
e7fKj+K3STK2w7oHsJU8rWfDjiIcNmEJ87/bGNwcB/3C3aBGuhagISvyI7uB7UMgIO4ni/o+kPBb
OFsvp2tF7E0tH/4vDSeOjgILQFyPluXmQfamaDKGkrASE7SgnCM64uzFYTXyMueNiIxTh688DyRv
FZEQkaIpp1OxBHIgq0liyOvr84ZxH6IYt+NKswEOtOuWIlZxzV9bKq5GUVMOgjHfbQ89mEK87cfc
Zg6Hj6xv5MdI7FbdDuBpTSQZvEdh4sD4r5rk2WSZzzHOMgquGlv3n6Sa+eIdVgWszOYgZctehhEq
hbtZ947LNNxrgit6a26n6SAJ3tnpeSmfqKUAOZA2eV+x/1idZfqWoTcRxp/U0fy7e9MIlJppqMbh
JydBgD2AN+f2/XUj6GsSPmmSFUfoc8jdQqv5guO1gX5Q+SLGfnG9cv/htnf0GQSK3VEPSPR0J7qW
Idj76NWxwSw6lnSYP2EilaUYgUjhJaG3smdd4I6DPYRTr70uxUzjkQRUr9l2zAV0Qt/s/oW6TT66
tXVWcGIihOBL0kMQos9XmcZ3dAS+GFIHg4HPxguHqQv75QaQrGO+S97emqKbGLSW7XO7C3LkdALH
K0Qckuzyy+7lLkAHKmhJB18Qmtr6jmPJhui5/I4D5u7JSvgLujeLQOyzbW/Cw0AVLolCKxwfbHEw
PC9A6UQcdHLUrvopURbEAvWRBTDV8W105WGXTm5ZCEO198wc+89AeUs7MwneYZAsdgbnb9jieo0q
Tuc/hfTlD+juCMDEGvWOYQPb3Ge0ILTynK58ruglEJmVpicwgb9RzUm7vQe1izmntNwEmlgA2h+D
x3Gn3+PAGTxIws7bAJi6oRZ1ja72OXVzqXagKrLQ5ZdAhahydHQbPO5EVWFvUk8I3W/f+8xIfTq7
C8CSHLledNmsbPjpbBcYim7V9cjYRJXWvPx9P3uh63v9/cgW9qVTAbuaTMA6nOswmkP1nyS4C6W9
29bBtSquNeKEB3FJl8Jlq4mg1SJya8JEXQL1ov2QD8fCHgabEjEGW2miAdmXSHHQfEDalm8QfuQE
BDWh2RMnI4gIuk3oTWAMVNg+PBKmjVF/dq3+UUb9Y9+/qwlJ0Gz7wUVYrWwlkSSKXpgAsXqAZaS7
DIOHFODvU4mnQwloOu4vXsaR3USiNrMwvXWOrIxBUC/C4KXt0MHY+jvmnmBUlXzCKe7s7VTLyxSC
V2WJ21FsnDEyuUpP1qFGJSiTqqiDfG9iPvZx7eyymKL9XS5OxkgF5Nfwtv9S9xT+avIB6l624tLV
zxvBv0qSftNFu40PpyRDLdBd9PXgM6pNvmg++B02H7C/sjWf3QErXLY7pbT6cTu1APKTpemzRKpU
pBMmcSrbjNKB+hntBIX4JSArxXNJmZqz1Lo7c5cm+rdhASGercSrgZEtcFZ4jeojf7px5CPnorpM
MXtMyMkmmYF8EcA/jBPmxnTEUhRd0mGz3KG1yl75/5ii/pEq2Wv8NFXVW1lptLNagwpv3bBmJIh8
M4iBy/iXPQFjeIQSsV//x8IadS2nrHhBeY/zNAs+9anal2lbh4wAHKyCep5gCZYkbteEXh8TvG56
hC9AY7qnukyEChn5QEz5RH86rtvdvIPkcQcVP5JM6IuqpxVBBZdZgvUhP0Lk11eBpPOcjiyEjVOo
VsOhM+fjULmXgr0HRoelmgKN6IWC4A8qM1muBeLa08iuklb+VZ59ySAsW9N5WTAqIMaZULtGoXJT
1kRzci7+lcvXAxp96bpmsU7UtBIxtjrx2N49bt4zQxlq9UUeIXffwqBWl33IUKZbf4sKsmyQXmXS
d2x5vEkFhXMazcwQz87bujnKlubKQNFBJCZtZz1mthspxouj4N/HhNBY7hEL3s7tWCs03Yxxds35
WaBEYu+KDMxtjx+6X6FYxLnbo1+Whz0Z/tsQXenZQO93Aktu4YQsEeXJUWXGoigWiOAA4CegDKEZ
/rZqtIK3SXHE4JNszlOY2IQJaQcZQqlPyxSkIg4345hI2/x4dUP8I4LIptrSo3kUu1VEaSKegr8q
akS/pw/VFNut/Dws2O9N4fg4rMCrjIUyJ6il9OgodN6M10pOGVh7/v2zKjTstVX1ucQixxFDc8/D
K0nMuS5AlYHgNmhp3DR9KlWxUFJ444ds++WRYK3PaI6ufjeOXCsVL56sVP+tX1kHiH/MONLZmQY2
0nl+yponjXiXV17liynFGlt0fAxrmM1OqvEqj+eTSLx4I8CR6fG19qqZIOUENgCdXVQWe0cHDpHa
6fzkzAmhIMHRnjkcCm9GxUBBzXKmDM5BKBY9ndnEixds9elkHg4vmHJYsF9mX9UKHXcZ62I0ppG5
X79QG0zlE6fD8oy4nrUjoil4VM7mGFNAfKEOD1ctd4c0Q5fWdHuts6Qdb2HZqbMF6fMHWIxGdaKr
76M03rLuwJOIVsp3Z41okqqcEtxc58ICDN1ZIQoUnHDxJuDhyvBvcKGRxXZiFu32K7WTzcvH9Gb7
32Z3GCgR06gzsurbXNlF3lxk+G72RukIt3fNojiohVx300nmU7MczeTJ4VozFgOCG2JrWxdHYhMm
/EmD5WCG3redFFkznnhjpQOMLV+t7+LHVqkXwfcC9G4y0CBALBnr9FuRVr0Y7i+SmP749UmaLnGu
wOpD/o8gdvFXGcf+IIupuVY/NgnRs/aeK+aTLZ2qGTdsBxBhJ1BJ02MgKD/RyYjXpPDuha5xK5lz
LLIxYUCml7uu8vFeMH8jMh2PpTXY2CFD1N/pX4XWdWQ+nujLaRc4Y8FWB6prUAJtPx+jR0F6/qvl
CYdHtjoPXbS7BstEvpoJOZt1aJLT5bC6H/5bjm6d+euXTICYivBwla6qh6xaH2a8LkXstga781dd
yTR74yjuKBJ2hj4bSoP2EHZnyu1mA2NzTYPqokz3GTtTUL/jkfjiTQ3y59dthF7KvKph0px0mriI
TYzw7G6Dc/LoYDnCGLo7WWOLmv5BAHdtWhCz7a/mrpKFy5UXwTPEzGPJC9/e+m1FoL0Gg3Up0CL3
DAwgvY39oCJJJn1k/kLsN/dW40CKS/JaXkmebHtRgAlS83p4BR+diV1ODepKNJjcMvaXF6cvVEr1
IyQWsi5mdy0JpTFjbpwbCPi05nDPReT3rYeOSl/zGGfzzPcHrgJfjVGQ4khrt0zLcgxb/2eN7k+c
VOJiClpFSwglKhECZRYUi7Th694mCxwM7ua+E1woCZ0ElU2ZSletKUUYaj998yqMfYtCijR6+6QZ
sWuEfvLCfetd0KK/fKT0EQ6tyHUzUoJsCl4zO1U0SG3gqDGGu+J5iybPAAhC7QAl05AY+Y5Raw8z
sB8Eqc2AfzUW+U0LU3Q3BrMM+14kwREq6UHyOyjuBE9Ooipscmtaf24K+BcuXfWriElYkiydmXzR
EMOCgy2ozBJhx/5x89YqxMraDwB7OoXBQteuXW4ekrrTVEDH9geqjD7hZXTjA4feYhZV11L0Q41c
5cWQQOi+jqHaVmwGqEp5mwgIu+czeeOCirDoCn1qFQ8HtrUENEWNqRDAi4qixjT+PUW2R2oyMMlW
7wDvCKljF9BZ1F+U9sfyclrFB4NQcIDM/FZ6fstBJuufuHQUrAg1lRoCWDYakKODFDzDjsDi5PvA
HigmvwjIHl2wlfN7DF4BDRSs06UvvhOJDqhBeEllceDGZm7dDpEwx8eLltA23r26oUe2AHO2exag
Zc1pT/2lSxykYUPhQrc78p9l2JE1uRDlKeVIfHVKriWnS6Ln5+ltChT80dL31maxeTxg5A59g8Gk
s3ImOhoSTay9ZAWDpMBoZffrRxBvmcqc65E0AfDuSjZkfhgW6f1EJjMKPZ+UCKSIP7wzpyIBQcLH
ZPY1RRQciBdT2qfrlz1RFMzO1ewmzHd926a8geueN0fLOzRlEPwjs7UnhacmduOcZPbFNXCPcVkI
YtRIIaDLKr86uFzGHGvRhmJ7673rbRUwI4iydpC32aAt+u4mfUzxesVmf/lt+2AeANktYLwWz/fD
Qd/cmSa5uVtyk8VWXTAyaqyOeIdU4e/6C7X7eggP4CxpxEofC3dr2mQl9XhLPNHEEmqWS1qHNWkd
LyeXiEhQRwuMGZ866OPePIMDyt0rF63wH8ScliqVG2lVXykaY6woqiMoYmGDH53jPL8igI+LMwuk
PUHb2Dysi8yoX4w6Bww4jigQGqKIswIJmcVjjmJJZD34J52NUu6JonUEqjzkg+owJFQQvhUepLvs
HxS9EebnUuArJESi2JgyQKVgg065D08JToUQ8QLBZUUD1SybMHGD9N1DMyqMMOBbOkZkZwp+Nj4T
ZRocO6oRjxmQNmoGOvmKCLuBHuOM0pb+PFt5PN3qz0HBksOtZuDV51rUdzBKufu5G3iiY1HX74lu
9BB9GktCwlAISE0IzBbxyv/JfQ//Ux77wnbaTCYuPi1+6HtB0zuHGQvQ9vxzz2v54QF9j8G0HC94
9nBCByLckylqfmr8q2G/YR+TYBy9eebQHK3wyVrMo39HXxuhf9tXvnj9fnQ6gggKZZ/EUznvHWdN
KHIRTsalcCHrSGD8E4Ed9HUtMC6tUZGiTQBRBJ7KM/sJ6PP/Rnp6Cg47vfqEcP9383np31EwrKif
7QpQMDSjbJhgCV0Uj8WHpdZ7+ORcHgWtltYkGPjvblSHt+R8dYkLaFd1Gb2GHDFhTPrzZG4gCj1Y
Z0vVO3gRT/G4pOu/1jSQHkFFKr+ZjF2Emz1m/B3UVL/Nx9aYdRduYVEX1JZgsAg6JYnSSbXWO0Bj
0XQlH/G2mHK4fDfpYMGVA9MymhaQ1mPB4+Ix7smQbt31n78jF2BeqgZP6Ol+w08RLEihY9zpXkDN
5tPrg37Jz6yTk03uyWtAB/SaYdJZxDZV9eWzvk5kz7ccQVzEhyb0OoR5ULsHIAO7LGaN2FIMWmw+
DF6c6kCuJp7AkDqlpDFmdpuxGNwPAr1MciLqblnxzpe1kuGJX6VQJeDcUp4jDI3GqnRbnDrVPC+h
QEZNZ12BUoDVuG7waYUoO0Bq7AMUXL2CaqZCqvlVpbF2Bu9XjAl6gP0T6dJW3ricM78q2IpyjSDK
apjJ4hMBIF0Yx9+xUT04b8YyzYYiY2erW1Y50X8a7dsNLQCo5loeECmo5fjoSOMOPCTKa6O7b8wC
xTDWFGOKzRyUFKZkeD8fHB+iBjxi4vmyOkO2E3PSC/S3BIySMg4c2GdEv71IbzJdRyc6JU7ndVC2
Wj+UAGckPD2Z3rHzuAUzrng9EsyKAVamdxLYEQf2u2qEkjPl0AxvC16HOGWYdopde2BkQ7llDcMQ
ZGHKvUEtfIvvMYDqjgZeQuMyKDhRnmdccjV5UDNTZKvWh57W3CB2RI87IyE7EDYN32xqmqwBAjec
a9I6wU19B+n28EttPG0YkdbxerFYWRkpmJOo/m4kkSqYeEdUVyawZJQQ5nmtsJ8P1X7kx/dY9WQN
B18QOd5GEqsgDZdTxM4fL7afjnPmrSzp6JMZwWbDoilqocGKenEHOAvFNwd6BbRqSxT0VGhARrzo
knAcvj7xyqe9ZHQwU/VmgeUEOAXmuWrUoWc81Tlabb0fQ7MmCByCXIiqP4j02wGQFWNtsze870qw
232zOYBfAJu7dpHS0ZlV+whFsUeu7yHpfLu8TVebXvtN2DiqRjb56WnA8H6GhCRLZtLxZR6SzScI
cR9sVOYUGMcIP41nwkNMAE1b9b1Q+AEjmREEKRqbrzZ1HyS1z9NraBpG7Tfh4/S+sjUjYOF0aL3w
kagvDv7o5RqZQqyatqvyvU8KROA0RBocNCz5RQcD8M4Tqyxso7EeFlrq0lcOJ0D9df6qjbZF6QWQ
Y8T2Jdc2DI+e02e9f7BL/2DU2YxtYOnQ9c/WG6/xZaeT7+M2jBxif2qhFwHqTkr+yXQzoUU4w0zA
+pH0zEI3yFBwUlz1mARSbB3S8mp5M9Ds9YlOJ9oxqZH59bYHxrjl3Xi+0jC7yUVKa1Vj6X0ZTCBg
EVZWVrdsRnvVP8n0vAWJ8JhNNskrBTwL64LVwBE2DdWQj+1mmpUmBEpFZmedjwIKIttUrk7NcqGS
cSdwSTLkMDSD91sTGb7JbDuTg1PxXpei1t4XQzz4OmqIoSaHv7PZeHVVdmU7y3O9B+fdvMc0G9uo
55kLtUfTWDOHYKofN5kah9Ke/8zVW9jyNUsI5KE2UeeKsVntApI5BjnOAI9mfkKCUC4aHkXLcmF1
pgrcCrBC/HSit7CxhpjI/BbrA/v6SgSFaX8yUDnfLVyqoLJD7HEe7kXT9ED1JpdV5ze9YH1xhnyc
6BRogQN9rQwtWan5Xt9mbqKyPG7cPrxbtRX/1ExUAz6ABCii65MLpWkLrMCDzeraxSuPUHYyL4kq
rhCT+ATA4NYzVHJeGnNcq5cOd8rpP81F+8znNt6Hh5SdUwF3Q5JRVIIQUOqC6jb6njQ6epimHXgm
UkGvXb3bW9uGFNny1PJ4a1j01DF/NHqU2QwJ39nlMyF3DhzFqOnlfkiouOwcbWbdVVzMSgHM/6nG
KEbu5eDVnt9OQYwR3JcEf1HhCXIQQ5WaJg4xY3BYqAdPcToCdpHSlp9K111NPuOY0GbJaNWiBM3/
aSaTM0AXuUr/mzSvyeu1ai1XdSYgsNYvtFsg0TiK9j2NYZc72aomZKQeZXaimfcwfl20xsrPa8pY
KnzJOVYM9A+R0ZyWN8Rl8asMRhJGCo3vtA2GvuNISd6GpPGhN9Z8NjRqWfhGyqFIMr0alFyibG9t
Y1Zk8l8DzMmqLwnBlP3KbP4xbvHVsQVktrgWjCLryVnX5O6o3KG/JqfuiReXBMVuaJCUSLnD0vGq
b+SP6RgK5sfaSKfxyM4Sk+c3k/L+WHpjR9KtmZGIjGkUIcjvGoZ34n2pmdgAAe0qSRFm5Q7gS8zW
jP+rW3+lA8RC1n/Gwu6+nIJNnUWKNsGj7kyvUHUFmLJOJWdTFiAaCGOuhgMhSpktoCPmlwYPTHrt
1FPmuWEadaF3wTvybx2ueqtSxf3ArM2nXdLMEzW2tCDu1YJEUGUZiJhk8SJYVmCgXBIUn04mNd+v
J0LdCVvsWOgVjvm3Ok/6bJyS21HlgH+NMoIamhPOTdkBEoeaoq69HotMfEGFc3YDTL/A18mQdHwB
mvfMw60ogSXPD/ot348spNoq+iTBkylQPUaRpuGXA8Qa3vb31bXDDk93h2luq/DF/tfkihfdkETm
MfM2PvJY6n/6tvg1fuhI/CIzGdFFrwGt+VoyOwoFJxLEJhd5S1382yo+uOXb/xX6EjKb6QE1fTYF
1kkA+Gf9YFzn8RGiCmj8/W1WtxFZiAz84aqW4JEwdeHunc0JQKGWXXhgLvor05HrRMyn6B/gaY7B
zavNXUPaeO9uAWcHSDwPhRv4L6QRdAKaQKzYGMxQZdGmLSSjIE+xLYuKRt40J1TjUzIEJCniuZ0I
/whcehYHL90dD35yYKvL4Ltsxp76tdG277Rh5GKU5rgnSakuw+KikbzggH3NyVcFuCb/97rQAtZd
MU/ylB7GivZssBiTgWtqv/BzWhBNcDQWN7UH2PRybaRBLlMUwV4YyZ2fiRU1zuwPvhOIQA5/ypBN
1m2ECco2AlMy+LcLTIjDt9rV8HWa0mhTWXSjra3CpKUooDte7i/mB3ErumMsdFMylskUvrDkxl6Y
Zun5+VTKY4WAyDh7hiQ+oRTj7+IJouZKcwIncqy93LW10z/W/MhUIF92XpE+oL/n8A9NU6/ofh0v
D6cwUeXxlpZX+cmzoVTbNOhkeoboSefBMi/tfTqETC5DR+FlQg2umcizfhLFnVIIONA6qjHOFx1Y
fZYyR5J4Lz+BJ/WU8yJWCeZsWf9EAq3ETAdRI1NqnGCBiBMHULBRvcuwmFv4S54l8I3G1nYMz/85
+X25LcOU3FDKGpv4JLvSlsQcu2/+D9L35jXqT80CSmay3Rp5DIQUz6HuiWFVIBCYeVxttrEcP7aB
ifjyj2zSpZC8BtIvfKGOOhl8yaCBP22EfCCAVL2R+UVJpyALG9Vji5md6neKnTbuO8lrDq8MO7lP
+tY/WmxoPu33hbTcBKuTCfCscYfuoaBrNflkG1abcJ3lHeLdI8GF3yk3PYpkARr7+G+Lz3of3szY
zkN9/W1YnMpO6bdmt1195qR1lIBkEl9OFU1XIBkjcp3BTZROfW4VIeqwxeQ68Mr9LMB/7yd3ZAkt
nJBU/El+Jql+sh76f71QHRwFjOOmFUVNboMNFDitDjaNhDUSw3YYZpcYAFVugOhPh1Fmc5jTG0Fl
TUFlb1VCF0TM5yAw79a/T7pmy3PHNj5apxaXffjJxk5Q1uVHppTQ+mFypYsVyXhtelYKAYoUQqVD
IlAd+ImbEDQOKAkr4gMr11QGMFJ95dkuzpNB1t9sOHl+TYsPE+lVTILB7Uv8puOpOEcW1Vgi16bm
tr/xx6SmMV2TkpkA1VsiX0HZVd3hvMJpc+eWrJbM5Cr8l9H6/XG+ZF8MBN14rpUeJFuHlMAQPRLH
18sFPiRANMqQTe5KwAWMLYYneyoOvxDUECD28ClYRS70h4lu5VUCc1D4OWAVV1+Dza+nX3gkBL17
MYAp6Q7IfrL5dZEdCJqF1WWpo3SPtKIogTx6+Ltt1RuxrmzLDW5ZtHGtui2sO2iQC0nzju7WAMtt
S6FrrP13Aj/fPC2B0E3C8Kjw3nj5Gal1pLYKHozlqZ5uLS2ER0iTylX/wRqj/E3aNRg7m6dfug8H
Q/PI0zQ+p54rZQZePcusub3ulpB//ogY0pn3UA2ZPf4cy1Gd6CwypkqXuyGIYiB9iScw1CODAyIP
ch7ppSELItDvQizgQGFJndV8/gvYnW7pQwDric8zinULrIj4e/F+4Q/6wUCtMLB5eGzZ4YXUZMzn
W9SEg6gLrzSh1SyYKeVz1mIiaIDWa8DUyoLIktYZ/YX3cLKthqpeF0HlkdktB+14rfzGSTMakNEj
Ep/xjAO0Qyg5x/Sa3IgZ1OCBWLrgRM5NpqMKQ+kVwD2dmDxp5M4nb55smnpoyi3ObuEsocpVHBQI
D/swbyXkZIR+uDaatr+g8F5SZkHxlULPvDq4Mdcsq+KaB5Kcc+0ggJ9I6YCg4dnzZjNMfRkMr2jT
OPrT2ZZomIPEhsbP01MXPoHUcM073N4+7OPLsHlidYySdbTqsD8Yl3E4kwcRetr6nfeJ1Ly+LSnz
uSE611mZziRwG4QVwom2qqrDTCXTYrSo8LDin9jo0xlwR4lL7dEffsjrnY7bx/j0SnDX90ekQitV
Ok9t/ZhxIgiLBYvdBpPabTriKX/MQh87/Hz+Q7aPitifegiScr6WfMC1aOhw7P9O4HOmGJicORe0
7hzpdOzJxZGLpjfMaaxVpW8Z2cnONOQLtHgZ6Ncp1/KhPyjg4xvgF2FPeY9QexcisghHLwNyhfk7
h8S1Des+4R8pRFDY3oZ9zoD7Ait3g8LFNuynxy2yOOHJCtBvUbeN8WWPmFYzxCbQ68z/gIAHoPdu
FcUBWGfIaiEX0UUBRMVz4EwP1avNA2gfazNIhv+OI9TDzeg6w5n2EokaS1Yzd0PAK2MW/lm5OGOt
wKnlm50sXwIVH03vwKh49dLKX2iCrK05eEREdggDwCYRYA1k0TxqJmkC9XUM1CvVTQ7u+etUAG3/
X8gYDaLmoqdTc9HJ3tSPovMTAApoa01QYXfrOePU1fUKRq3eQSkbFYOCmne7KtwTkA+Gqw2SonsR
Z9Gfaj6akAqdj/XSFLyLKIdYYfASxgT/Iuvlgl9Pzeo3FEQfgdKD2buHoHmmqzD6nXxKLDZFL3tW
k6lmJNU1xaML8EbG2V4FDIKnt/76/r9u+UoW2DkmXQm77NIrfZwLnVg9R1w7j+MFn0YLei05Tuq4
GdgDjq2jBTup+Zs4uNBzXZaeb2RazDLcXgCXFv/2Vd2o8nN2wVleK13RANrGER9RXegzNOg+DQgP
TXgjpnS47kUAFmzDpuIDJTdslbaKWcNBMmDA72357tD9H2TeLwxc2m89HvJPXX4J/I+460knEYzo
vAJo/zaMY8gE3XOH4AhpjdRDycM9p4PAzkTp6ZPkcvVm2R0V8DnmKt4IfZ5BcPZZX0yqfdqY7EZ0
PE6jq6nxyXq8ndm5DIsGPUMx1llyVqUMRTQMBq6JR5Ytg9n6M5BB1heygAldMML4ENs4QdGe6W/i
+8y/afOZdtPeOcQbX+tRxZW9IQ+KtZe7kbNzK/hs9s56ppO5lTDPE4Q2Jz28B0Ryy61OnOwQJCdD
Kgh/ntmV02FfpsFAV2vkuMkygLsOsaKqeemmbtpUO2g4N85mEH6tPFSgBMRTKjVCpomkE0jm7QDz
nZAUoU7tkz/lED2QA10fEH1vbfk4D4PUzibRUmZqUU2jU0v7lBLdtY8wOstlFFGZEClCAk5nKOfJ
QH9zI+lAHIHx5Lii3twQuBr/VNFJZ2gHFiBcm1kkJM7I7eS1YZ1Zzt5iHXAvadLWmLR5SXq+17C8
tragXomfL9+VXk9TlcQsSUSG88gBL2iZnbYaxTHWYGx4g2YMzoxmD1sk1J9gOhCP6AVDEF7wvFAS
ilbT82FiMA9TJ8tqgLCvx6ghOVp37e7MSc3DMweYkT1BBD3+Tj5Nx7fFeal+qFi4gpoU6Ru6+WV5
8g5fvOc2iehveL6xXoSohI3UC27BUe4NEb48AgDLw1CmVcs543/Qwg1hbWSJMOKVanC9IdzQnkvH
cqJD04PzLWMN7Xqpw/gRucf8Brez3wzivGgkEU++QlQ4RpPi3k9bZgAs0aDCh1VfT6BOY3abHUzM
8aK4b+cetUJR4qA3XWRMI5gKsIeiLRq/Pkrr54EniVQS/73lIs4CAoHDek4/EpWvK0JZgipYAQj2
V3se7U9N0Pj7ELRXH0JNRej+178VHmKFFOs2ab4x4jtgoW7naaln5npoCzygMDR2YpNLTpeXO3tj
GyLew0WkgptLIju/ey3RvuoGgy9eHTrt5geFjP5Tv0isX/khJC0s1ITS++wMusoVmUAUnajkVxr4
bwjWPp5u26G7Us3fvvE8iwRe4/2/9KlqRLApxVDGn04f5EnIIsfFLn7gr4CeW9VOHAwGWw3Pojos
WNAYkJRQalZqDCWqngkUt8q8Y8SUjlLEoSfkCM92SaefuwqM0Jup5Vl2JKMUEELUIkimz0xGKjtF
YoEV/Z69FcZXu+6NL/ZY4IfOGp1geVsUD1wQmbtrZ83XduDKL/pNuKZqBHGquoNoCAVLb88I/+kt
+Fh96ASN2wp37q0Uu9OE9S4piP1yfS0UVE86gj8Cprmbe5rs6PsFmb8HRaGhj1rITii5fehHWpyW
sUgOeGtZkLaKGh1K6pMG6/Byf4cKcxLROy4uXge2QrymKDvGF1OjFS3e9Qq69+UHJq0EUPpoTobe
arVQAa62bZJw9dlnI7Eg5Xvjs2lmGSpPRW9TiH7VkAQ1W2uMBhHf5jucpdrKy0Qr99L8alqCsYQA
2O+AvuWzP/X5K9nFl703LyhKRnTWYBJvnXvs7Jqkn2kUBP4ynNlA0sU/x9rYLXf+bqRRPv2RcCyC
uqptFEHsM0Rw9v7CAkFPxQyeSh0BTMqV5ewCW6zp001IdNhp8JpVLklUGw4omcbdI1sre80xrI8z
qFDVhPIOSmHOM3M7GRwD8RVss6T/t0GfI9u5xyoFX3k6xFQDXVvsfsb2KGtcMLn16n1G+GzSpOzs
myetHAvxIgk+R3J2Al532ojEYj6X98WUoMs2uVcLnrWKvNuM7K/BbuQ5PxT8sHY/qQ/hc06mSnE9
a4Su6Ez+1ahHfV9hQh1YH5qJQJE44bjdQn7Pnm0FPq63nhiBgsgvem9qmy2eiqcrBKCyyg6mplYB
KDFhTK1GInqnqcE6GHTABxNxBuc2i8O2XQ4V8q9NTlKlTtP47h5Gg1GuNCsbV9124y1Tfeh5laCT
xkjeRZim3R5Gpv8SIlZjheR5Xj3mMndag4UWq2NDesN4trseXe7VYroJVhQebBbYzNsxaT+KemNW
HJ/foKgVo1bu9cV+yvMT9C/K/8l/Ys1UYni/YmvgohpLSppKUhakwvfcPxZU/NSMO+jTIl5xWTcR
t/9Z5+Pyng+4rFd1qACSWQqvzHKDYfwaf3hm6r7Gk02iUGs+1o2aGJm6IhqZjTFcK9jjQXPajekz
1Hw/UVfxoTfjbxkPbcQF857p59lohE3gL/6BjdJF/x0YN4ipKORybspHXan8lu1tLj/nJmHa5XVW
mCCkdP0Kd93PrdDS+UgamHUeJX4AT7n3Gcmpxa10ZU/S1DozIyPxNUPPFNGtIMfjnIjZDPgHERpu
2Va64la9tF+hf1FBn69QuKrUd9WQC7c0R7yc556pR1/ev2PGZYySy2pMFQr+PVpjASnHi59B9s9A
VMDpzG+kf4bzQTQfwItWkonESCXN6T2TWOzn42qCPLAI9AqKx6P+sRafJ7npG5FJxjZt7tsJDV/3
QMCAIPMcDgNRr+fzWMTBynoM7KPvz2+1wTETTp3qkKYuw78JXTH6Swrqu3k9POFU1UL/8RLaMdUp
20UXieNhCGZYvyWMGBawvIh/23DhC6Xqrilhnd/UQr3rATwuHl/NwXIrdlBMJbJFlWSkpljM7Jin
EtzB53rHImpFRkMzwfwb4jcYcV1r2/qZ9oEvCGtwNEXj7Cny7gC+URN6n/suZQy341BQ9C9OrpMF
+xDWNmErIT3JicqnhNiYX+2kUDaGa0MMOGOeGyVjylpTodx2V3d+ysN9L3R8bqCvSuuhJmdtgxXu
fdVUpVuVWI0vgxcLxDI+MMvAeiSSnAD6QWf4HLHN5sskxQhoKkQobGt8oIPwcvWTrDIYLp3fKU4B
W50Iio6Crf86wJ2Tzw+9z4TXmxf9XHyNAaeUO4BxECpez2AzYOHEFj1zH9UiVRNDGwl3qdo6GB30
bLqiIpiGiJ/XWnSYHrRUh+C9zDHpoCu4MUWdvwONpNX2EPsezvLJXV+WoqVUhMrC0DiD2CxmGXwh
J5MdXhMuNEQH3RCeIu+VOfMKgwf2JDIV8/uu1FMgzp9Z2lf4ElOhujHhd1fDmX30gQEnwEu0X0Ez
LjzZ3IEVR+qVk5VLazYS9bAhDAZCrOt29bHYMjGbHE33BToGxbkqGUhoPhqK0MaHo0B827/rOzpc
UAqkv9GviBV/gLNOG4XWAXf2wwMXe9dl1LlgAcmLQZev+0jdW+zKR2jZky9Z+3NprNp0ktunxjTn
odCWmDw4tiy81YCkF7tmhNqLAzetxRj0uxdVOOH9dU9m6lymvM7Igw+OIn6FSOb11wBlKQ5ddXTj
wMfaMOl9ZKtI93R1bKC2wVJUzesID1fIG6sYSGFg0myZ1rM+BnRpJYN/B5Fd4YX+JkbaC5FeuhE+
Q1U7spuzXup+XbUCBuVcJ9qg648MDuP8zH8Lf+e0ZOdtpJOyzPetpb+6AnHHKCemis2Zu2f6GQyH
lCK49Ee6YKuWt5QSd2ZmsP84VLuJRM2B7thRZFuSV7I5WgxQbI0Vvz8w/I4h0cikiv9YdnC3XKvW
ppFUIogAfmOjtrytFsmMN1Ojl2o+1UOzJ5N0I4r5si2SK/r8UYcIVRG33xd9j55wwWB/Hb+491F1
CU9WWzLzQAkES2rCNiHv5QiqlyzWz2FHHe8PkIJmYBzcxVVDrOmShaqmeYD/oT+bbqrpkhXDefoD
fkLDDaRRAzDfhXF8PLP2gq9CI6gen42EaeeNNzHQ4wKlNt2bejiwRXPJL6aKDO5spC80jcmBHJGb
SOITp/Jx7+SC/OQe+UZ0bDbjoqCqglGgpSb66a8e94v/5pG3y+EiSOIWmhUU37ysadqufXnQS1JL
WUQ+XJzknJdsbN2HrD0lUrSz4YInH3tRTCHI0g0joYw26/Psnchds+3h/8q10cwdYxKTNz/wuw+U
xVFoYUIJQJi63rt9rMXLtdV168249TfRsTxrc7lxlHwULlN2TW0omQVW/EXwBQ16GRrOD7h83PFI
GRMeJCQ3Ltesk+CocMB0QcL0TPcyutRu+EgLWJ5fhXT+ZtOPgXRgnSSCzvmnPV1AmTRAqgkufQaz
ontVyKe2Wi1aeRqUX7xGrZSib6q7pKZkYxd558BaWxAvYHH7S3KTMvj16ZIuEeR8cg/yVZa3eXp+
bskqHel6itMNLd1N8w8GDzIwvtHy+loq7KfXcPnw0fyYAfbWRzfvVbQjcISTmV4BffaA5kyNZosJ
aujxzE42cSigT26YpBF9eNlLBGMu98RZqZRtjxz3DSTRj6XvPw3LtshH2+f5ZD553rJ2qf1exU8p
6dh+csMiXGiia8xuQQQRuQd2mIwOGfTgNr6FbCpvjx4Dzev96+QKA/WfUdalzgNdw257MMU8MxKQ
ZhMIcmTAAPBuXHFno0kKsB7nKLKzm6Te/+jOCGlxkHpYsg/XgDdaUnpU+1epkCYpIaiH81IWw38A
m7OKOqeLTFlkDm+W6lX3c7wzJZvoIMAg9H5hD3h0Nv6kA2/5cpC/q9HJFgVYxbo3630spKeNJDYG
eqzzdApJ4yRlnK4n6S1MpAjH3Qwzz8sFSzbM0k7fNOp7sU8sL2riFMaFaHSmszLk/YTri7eo1vDI
ptsDrpcj1nBBLxg5q86qtCYe25rxltNO279S8oUqlNVA1QYmhphLtmhjjzP1qwLYGqlKpIz1C8tB
CuDRM9h31AXV4RKfa1I2KpyPCuwwJe8QhUSG883Icc6EoxvkAWkMZkhqJaxLdSso31AJFRNcDH0p
7M7zusd9bOP2x1TAi9YnQZy20LxnLNq7tNuwhmIc1BPYDs8D6nhRxNmLz6JTk10MwkdkYbc1AvU+
oL+xGbKvT2IFL1E+EI9udzT4uZ0p22r3pWT+EkGg2dx0MSVf0lt5Di5k+34PN2GtWNoCiPOi4LLN
cC0AqIyLB9tksLyk9hh12WVSGM0wf5BTvj6FJGyIvwdukoAPC8KsvTUplkugwonR8qOoTRKTsrqi
ArMEPnZxBq9qVzcZa7lUxV6sxvjUNM6LzDR5fNXMLBoIno5I7Nvk1/PgFhe3F6h6zYeLB/Hh9lK3
/mlRaBstWx9PqnCslbU/jktiYRwDdzHXhWmnW8RieEWXvDe2VwjI423L6t5F1peA3cGAVfbb6ZIp
3InHP9OQ/UWW7KCnKFlR4AOUPcWP5e5vAL68vvSqJEFGhkVIs7ireTlsG7MsIrO3wp/cl131VGWk
R67V30oBODXFuAu8/DN2idc8y1lvs87r4eV9gcDa4wMJj2ir5tEFRzwCvA7GB4tXFVjH8+lYFLzg
7FjTTTp5ujUvVXIaAUMRv2FVy5CkrwF7zntZeVCYAw1VPFfk5uv5Fy4TJZlllS/bv+g+66zzppSC
D+cBo4FHLMtHskvw0ZEECPvl0Jxkqg2rVtqgrZxwwn96RGrjOZ+JqV6VruI4tAhrz7jON+nLZhL9
YdPPpsQp1yQ/ZC2TSnF56fOal91qhRH2MHZv7UA9NdWJuRUe+Hl0JDQb0jqYCiqiiVfqVbO6ficO
aEr5GE+OEG3AMsE5PaALCH50O2zlNVFYqNljW6bnPYV2OfeHf8txAOmsiCNBK4Dpbffdt5VvR6WL
EDgKDWzBCKlccGIl+xwAfpmqjAtxvdkPmIdtfJ5VkDXML1s1Rw7ybHPvr3UKffGqWR4LTLEZTAAn
c2e52Nsn7WEU/7DZrkxGrHgSNP6htscDGkab45upnZLNB0NR+M5Tfa4NROCU9wJd04jn31LZIBCw
t36ialSGwPOuXAmW8Jok1oLJUki71B2TPE5gIqdMRXR+voX34XQTtXnNxxFuSeXf2VZ7uA7FzJag
znsVT8UFVUbrqAUoybizVA8FHGin2lseweod2ZxVSORpEkZwRyV+BtMb//S8E6NNF/L3zkCIXsz/
mQuHQ3bWS0PVtITJFG7mstdouHBSaTDyj/xH+2ix3cFVhMPJOiccrgh2RdadOIgy3DdMdLmIMlEd
JT/M7a3DnOaTsElypHn1uozzvz272pnlstUjHC5BRLSzu6M9oIDFGO3tGiA7IO4aQA0qY29qJR36
eER8UVutZBiNULi/Ogcwlwt3MM2MVI3L5hhnRIpQhbu1bxX/DYGLxb5pRl3B/60uFmCikxho+XRz
/UHF2/+u6I5vIY74W+xThyNudTtM5tZjaHi4Jz0WAmR7AhUOPMU9N+bZvP4+SHM/CR9CRavmfJpD
msZ4ZEBo8TA3tB5Nq1pNMQc8hr3Vs8QCCvCVBEsGm+nPPDMXpyhN/c/fmgKv8pQYt9UT57lyg+rD
ndA99GrpCUacAs9m+1I0HeQhsT9F5JbwQVtHbdtyvYMSKPubwzFT6gKzjcPkgJaF8+N/EKT8falz
pfaBU/QPvaECx53IbbVtHwWmPuEL/n6pOqx/VxBPDsbSCovGgffHoqv1RulJoqjYpy/8PBC4beWd
0afxrVX1WL2+0ylwUR+A4kK1Je9kcMEKFMShBQKcuz3WjFaR1gUmw1pxkIGxi3qJzl2uPSrPxrzY
ZSJCnYNYCedtxd3FLTKfonxXSJkSnhPh5V/ngLtvPWfAN4uIUoYFASMm02Jt+QFlVOpHiklWv9i0
OBMNjT1wvqcGxvqIK1yo2tNHtqw+Ojy8+GWK1O5L/8IkMWSFS7bYsns17PvhkxrBtSfyq2DjYbO1
ZYcgBxSruRruhhXPwYCpwWVXBmdLiH53p4tHFZPY3XsEPDVgzlVL1EVwo5d3ThUE4fYCvljDrrWk
sqOHsIc/rzW2kfAgBYcgCFOqp0vnpan32Qa9ygYJDdwtGuvHUhFabaACDQog/LNQg66kqnBEeqS6
OlbcJP2Y9jcapXBQ1YJ75eeeQJSbohidz6tcj7XX+zg1aRUGraRnF43ktPpdimbrGETr+TH78rAS
56P0ByTailiX/nKNKNu7oR6i60IpHxnzlyqZGR/Jf3Tp7Bkiif7fA7j/ipl1e7hTQfnYEJFNfO3r
RCBMRcyaTKebQ5VWQ+IVLxmGvpXgIQsvDSERs2zSRwpktIhxUygV9OLpM+cHCBqj7c1EPEAtBTJk
P9BlFU+ZPvu+XDeaPrAmPQ6Y/5qddy6kvJvl+rA3vC4s1CE5uSbTDraMKgytlnhvTpttSdQ8z6gq
wcOVvV6NshAbmdNbnSEwAphPdDkaOxq0sG40QNEYCbIwrT3QSM3H7A01qLZu0GbVVa1w7bTy1Dmb
WSKKXOxTPvcQQq0h3EF9fcZa1Oo26ztq5U4j4/0ZeFJmHrpTJXEwLoCCd6UzcF+GrtmyC0pNOhFt
YZIZ5mg57mI1QrNLkf5HsboHyS08qvHNjsTjtc/h7lywrExVhle50laq0KWPRKR1lTb1/aLv2jdX
ysfGDWsDTU/2x5CMltZxl8yZ4BUlYuSPixvzY8pwHGa1ZDlUt+Fv8EESacpZA3xF0xhBrj0JgzrS
uEOnrsiqPPhCONmd1hN2vQHkpzvOvuhcArZDwlwaPHuiktniGlurWNWFkRoALRXRn8hgVds/Mi/t
W/IZHOAh2h1b4S4FlhQqmBR47nD20IAPy7xINcifQF5IXl5mWSBRtvOkqnVuacSxXmfuNX0qVtlC
ALnJgx/uHUzM4hZnpZvR4bb9Pboj7eY5usjMx2HHNZu7FNFA7am3xwD6tNK2dxAAycd/kGyCwJoW
f2a3wQ907BiSHXvsgea1PAvml1wBD1VN9LzVmLxOvvzk0KV6cUnxQxJjF6uiOYx31h6ccRoIltHe
mqIhSvz0DGmaZtiEJX6wbspJEN7n9cqUZ47txwyuj/F/DhV3gN44f3q2p3+FBRBSB+0Cit/+Dou3
9Qb2OXi4ICW1Spm3BAzp0UB8g51YC0Fgyqj6ToYHTiPATHKcVF2vv38N1WD8s/p6XJUxtapk7gKu
F6X681uf91IQ8inY94ecm/soO/0JFjYCx64y2X3E/ytwZQgfsEkH6w4dO83ncoaXmeg6BnnZ6cIK
T55VsCJWY9HC3zcrv9/Vz7y8t6dzOAKkqHwniEnPj32SKv805CmboUoWgvXap0tYk1RXU8hpwEpM
m5a8/YkTIfxSxfukFSUv2ws+2mjE+ORNnmdGri/42+xWu2/Zu59VIvSRQ/6Ft7cGNDTfGap+2IBU
aCr74tGw/zFVb1VOwhLcLVcec0PZ41qu2vW7ZKb8adq8GjVt/ZaenmfKmsXxLzX1R2AzlDPskMJY
OakRr248QTrjsFRYkbffQOji7vKvqz5SBOCnDu7reT5icpsFgy+Ukp0RA2d/fuZQBK6/ox1WYmJA
4PUkI5SRK/K7NQiKKMjirOx8FYtTfKjfc/KrFGXWt8fWVEWKfAvkE1/zuIMP/0LwcNWrr7fUqGsr
L6ABvZAZeR9Y3QBJOwkhfb/KFvVLfyK0dTuItXbJLSvkw4KRbWh8nC+XyBM7Xku8q2HzqwIuIRde
9uQgqTvNi0vM14S1TVnrjsMOsjh7U/XGhnQAFi3IiL+ugT1gyDt97yf/hTjm500vCEF6OXRweM2l
XCyR9aK1BuYLD85Ho8y+EISJJoaIXnq+Lap8uuf4Fdj5MMpDEg9ra52E8REIVlwECGMMrH6X9pXZ
WWoQyY7gVCqpTiPdFFPXGbFxIk0LhcPBnHFq8ltMz4Tw3qUTIvwMljCWXcLzr739Hz8Bc6w76/AD
N77kn8YH87VDgEBcxL3lIr1np1RhAhtNBGW1Nxzpqcrk/E3qUG3TRzeC0HCVGiKZOOKI6W2Foo2M
mCGfTUpj/WOIKuXS2hoWIhnxtWkjokthUAXXVB9w+Ir/dmbtspTivPz4TK7b3cHVok4ngUQpWStR
CYUYSQRIsetSMq8Qwrf0QY17oeslAvP/dx3tInNy7ZknsE8KXr+LGD70qDmxFE7lgZVQyLGnK3Sn
EAmzz6zF1GgV0DAerXifdpoP2I98vB3c6bpZAL/UwDjIvS33ee/C+mUHZ5aydEjezEO5wzWmwTay
6claaima2oSZ3E3yAWBYKy8/Fbc0+eafHeb6MmZo37xqC8R126AdpL25jD22u/yb6QsRKBeDD1AQ
nlYtFk0j/mvT0uj3sWuVGMQY5HUF3kxZfcmq2957ZggRRyd5AK378d6G8DpPvlQCTSQpQPzTJKU4
RS8qz00u/Q4+4mHmkS2ZCF/6uYod2kIS1dz8W4Uc4Zm/jGdAvHm7wCQ4moImZ0Ybl7ydbx0J/nOd
38yPaTXqya7GYeYz6G7i3osuf2uJLYRuBJO3ysN+VN+KvP/jE7Ubx3uEn4lPqRKr0+iUMil2pX4B
pg/rEiEa34pTk2kTmz++dPR1P6j5SBHHg5KzabAnL/aGluEHoMCmlsJba7VP4xDhBoZi4EZiwOaD
9modTLtHwY103oxdTYk2hnGaGGsLDisdNdImmQHJNCMp/pLFJfqv184xJ3Y/2NE2VMLa3ADxqLx8
25sTkzPAY+qH+kKKaOrfQCfsAz4UY1mTS15aDSh0dbIMoIb6MrVn+OGaYWxoGcawYU5idNe7lCx9
ovNyDD+7wKaRF7WSyNn8rfiWlA6Y/UtR5Dt0vJBIGDgrsKEKwxut5EXrDLiocFh4uihfYgyySqQB
i8Ia3Hi4WrM5/67CA6Qva+8GePeDKTNcB/IbmZowRLff4xmEUCHCoSb/4MYeQ7Q78Ur0QJ0D5lMW
dlYYGXpVd7SnQVYXR4iYQk8oDq31YcCGWhcQcCThEHdLiyT7HPZ9uaR0y6A+lFWXYk4ZvTsM8j8b
EQwhL/Wft5b3urhPeNHmNo2R5Hz8UkiEHnrA6d1chttfTJM4WdQgZXo3dKt/axcA40HVapMEM+E4
iRaID4Gjs/ykcQELEumhz18TsrEUvv6fAmTE55HJg0TYv4OZDdppfbV96MOY82+s90CIEYNJlmom
hfC9OpRzJaxz1uZT/kiXQEAJ8r5AhF/V92/vNA5ZrqydBOdN1oYS4GdNAGWR25BGW1kXTyIpstPU
J1e/Ha8HPU5JPnrR5RgaPd9X2QuexPvUL2aM/JWgCQk+Bs6OpvVTFYQgzJuhZ7k0FpRg2cu3WYxb
YS3AOrD5OfoNwjuTvVIJXj4k0yF8HAadwW00fKj26eJyCdYyn2T3w3bMphzeArHgrsMQMqNky96P
UtdGnZw6YC2pMB08zQr4yew0cRh1A9i3TEmqC0qab4dLjo+2kXMep+w4ixX1Q1+N/IgjB1X+itbr
48i7t0a1PmTgbdIa1sl7GRZDlOAX1qpBBlaRnGTe3HgXUi3w8ZLe1ZzonFc0NVEL8YbO29VjIbyA
LIdwLch10CYYu7HUp0FlGBo978boppmfsNA/7Vh7KSdgkV3HpvUJ5vwrCRun1VyHv5PcUWn7WqZh
XwQpSnIi/TdfAufiwEplsTkxaXQ0ZLqRdJ4GivUqCi8RU1JXWwBgr/73ZC9CroCliLfSZ4P1xME7
o94z+mqpm2w3lwaJNMGhL8BhFk2Qp1b2gaAq51qDRXwoGO6eP+aaqYi5YQVvjbkfrUUHfMUTXoyZ
Qez8evwVkLwk2yzsiDatZ/Ki5esxLSIMcoMKE3jkINsDJNlk5Pnl2SfNsJApQAT8HKfRh9ADboD8
q0NFbuICrDaWHVJIGYsSFu864Z2kAkT0RXHNz8r90IIY3eGFxk6bqB+bXSS03pzzEJe7rnezFSfC
nrD66sCSniqn90pvg1fTiHT0Q67lgh6r2LYxyOxS9OGtq8HiKIAGK2XrlU4u5Dqxu04deRNfaXif
5LNfeYutuLITky7JrwccMLFghk241CJea5jGyWnBRs+WZpJnj3ahjV87Gx+x1oY8zB+VYSZPaW2i
vzKQalqNetcAruDendpbD6CziAt2M/V525UtsjRv2/SL5PUjB6uF0k5Lgug1cdCIwiZP8gsKRnnW
mU9MfFk2uc3MxebgWZyrF3PtJUU2ukYySh/T7Dj9i+qzbgzfuAkLN/npXBEM2CTbGWKmCTcYr5Cd
Ipk5C+LWSXXKBP6TXq/3YTfosn6sOWHTxlZ6JtgVJ06NFACfLokKbXFW7PzjxEr645DcdfI7g1jj
KL/PMOPWfthJYiJ/wohoS889oy1Xjt3+1ky+NCnxmMEgTnAod/3ySSJ2rZxbmt23uaJMBwfR4zQ8
56t3B1YVHXPUYthN96nRESDtt3pm3FmiU99nVCD6EyHvgzhI3ho172qhuJ194zgMOTKmtsDZ/DsK
pda6qCC8nN+Dj+mbPJYGjBbFzZnThT8DKeWWyjkfNw9Ffxhbq+wBcinB1wzpnfWKu6sQXi4kFEfT
6VH95/eMgkLdBmPvHKRdIP5kTkxaz7aYoSpjO7hBvI3JZg4nfCLRZ8JCwxYAeGKosY37ShF4klKF
U22YtzucB2qRIv47U8Ocf98dNwiYL/4V5BoCjEGtWCJIHT/BJpkeHCk8OFa9JHz4K+vpc6COSzfc
NZuymJE0FzDJ4n/b9p7zsfhCTqTxKSJEABVSvF316dTPqJxfE9IZ1iC/4amGbVyKhBnbucgMbNt3
FN9vCsFcAgJrJmXX6Jk2FcOmLbAqr/Er4moGXFopdmgQQDGTfzlIFCwpPS+zydN5dlH+0Ni5H04N
s81t0Uyml9mj4jO8QYFMHz/ctznUMcXuBcpsCEfAzn1eQQOcOeUsGY9sK07sXbf3Z3iJJWxxGLVq
feHvlk+GvU0sQE31yx8urICS/BTNBR2Yc7TotVmGwkIs2DscTxnaPD7/guJ9aOeoMyqOZ/LitPEj
aL7Lg64bDvjpZZS4xxT+CHt//udmCI06fvXjlrPoVhUEdVRwqixib48dPWdLSmMv0/FdF9rIoP4j
QRYdNxmKGkoSAGd9Z0HBfFmnPOoT6ZUt0Ko1cXhnfeeHCpTHaAkeh0ADLbtP3Z+3P6ZUQDiLlJBL
VQSOvh36wbCdUihV2L2cp+4txAL3BhRmNvfNXnvdg6BTgrEZJX+lfvRWV1XIjVHlyRqAJPbfya7z
gGVZYQG86ILJmTfU4o5baIzb79J7fEovPpNfQVny07dxgAzIjbhJXebicX+XKjiiusM4AQ2S5Sjs
ZmLMX+3TWnGt8DjnBDxxSzbn+sJpXLWczm27xZBHwWI6utg+AQbTbzRPOyh2eU6/iKgzlPnUnxQi
DMxQ+hldwsDUFiFgxJqKIUM0je5hV4ZTlL0dXFOjnahRRN9oIG2071+V69gcHZV7kNQduFLGCZqs
L6nxMUNSWfo6+lg6XaxsSUG9eT2mAoKyaBx4+SncCbwAt0s2mI2cFmovCcThiOZxoBiL3gD099M3
ySokWC6qnISXILQGmLWWH3ftf08C6dyxWK/wv+sk+N0PiGc1I1EBk1RAzl1rOPcDrm0OtHfcbDiY
F7j6a2u7nkH0Y7SroQ+OhiUeYVTYCdla3PhGXNN8e5vPNnoFxBoLYzcw8xLrdInI2r5m1K2ia3jM
Th/4jJk7XZHZNIiYZHDaG0HU/f1r/wWFReXB+dcHIKf3U2zzWFlhczAqlYU9s8xv7Lyai7aWrDtW
1niiATUba9FZbvqLHX4GBtUSv5QBiupEmtoi4XQtJbjGMpe3tpoyRVcZSQfdQjJaP4WDQo3HCUQY
sJHRiZvgnFR5nWcPrnIEyNbeo2NwpqOaexlBZPoE6L9ieYSKwuIX1WMdMeYFd1gf5zAEnWcpontm
dToNIEbioDbz/TD1IuQCM5W+kzjxYaLl7TTHn6bq7w8g1T8rGFG8RdNCc246BMLLFueT3mYCVfGC
21zgmCi6rRSEG4rm3bRlSgX8NIxWPlY94Rd67MuGO5BsN/nnECJ0oxHl09JhCqnOyvtlEk7JdqM1
evIHbPkxS51skat3bmJmbwg0Nm70vO68Fl4C2jkKaQcvyUQgQu7OJtlg2OVdiN/DXc6HUz7HlWZK
8esLneAqLWEpTV4qiD/rZ+mGcSBtPmn+9kIO/qc6nYO+r8CIYRMJtDVZCf4TJ6P3RkSxOL18Mqn7
9ECf2UsxJw83BVxkMvjPxDWtD17yB++0hqskKRO7SV5LIICIKYTv87hvwxVe5zM/wdyemB8ZhNuC
huwe+zPxnW/hXHHee3WD6FwMZSHO6yZvDjPteHkDM3DjNyQEu13DIYLlNUhlP3pDey+XRxkECrYU
RjPcEwJPToVc3vYTDgFch9xBM/0UGEzc9eNTdVMLDrCtPrlUvti0H+Bz1ZIMI+c3Exbb5owYiGUy
6yp7ZPERTCqhO0+bzJhQuML4Q+cGsSA5TRkun6YkL7GaX8zdgn3BqFpLDZj9865D9hvSFUgoIC80
CjHOemdlWM9opYiNAGBpk+HMY8QLEJFzcxy3CNCDqqvKFaOQ2lP9Yu6dv5s7IROAHEgmbfX+Q5r2
gXHpGRZ25uAgDxkx6eVE4ltAfreqJDre4h4ZCVP50AZUAP0A9Fjawbv/J2WYLXhL/k1rgTShcO/M
lG0ZD/FSgcveN2hsdhYWC3fP4Gvi3ZglYwm0cuxZOdVTdSUys7yK2reAGpgL2t9fj35yADLP+vrw
3b5f+mo0MAfapbRJlvQe3eNusiwdKyhVLPKikmMJWlqYz4MXGIKUzwkBtZZX13J/A+jOE+TfeNBb
ay6FXpw57robFQXq7ZMHgx3mHooBS7I6GkKoLT2hQPKSS/MFsdx1k9kS7xD/MOU+REjz1CLmAJbA
qIZpS1W/j5w/8UQbmO/+dAyMyXOm84DIif1+ArjysW/jyXBRX0+tC5x37iAtaGFKbWXWI3xQy7Sm
4Ex7s3f4NR+VuauT/MpSiElrUMdfHp0CxM/P8Rh4mz5TqhzmLV1AzwLVPbKtfPnnHYTtLS3gr0wq
20/i4mH1gUUCZLjG56x94ffQcjDa/ZFuFywci6TP5+OK9m6hePfmvNNUuazzrceFBzAVdZQ7MNvF
SyBIsyCvp7W4jUIOkGZJUnyrNUU3DUawLYHVLqFk4XoAN4jNAUUL/a8h3WMaNGGNDfIHQ9WvzDI/
3KsENOcX6LXhU38G03OooTNhdJQr4n8vL7opzq7iefRGqX/UBMkZXiWF7yhns62hq+RJ9ZPChBQp
uqHbsucPOatUFy3H3/+1FOBrmJVvZcT3gtEvyEIjMJNfF70d1BEnORoa+4sFMnABFaHAfzT/FW5G
7Sur/gwUha4zfqNb9UumeNEZLO/sSfvjWbbIG5WP1lHi5/DdVx8WYtbzXVW2v1jvhEkDpAJ611Ry
D87qfMvufGnJREmOX+e2ph7VYXNRue/sXlFr77XXwocGfwTpkMlvEZzst8bZEo+VMRrmwIZGX5Ku
pFH9Rv8NcAnl7deTDtuQC5DSM+L+qjFrp+ZpvL7Tn7yDegPkq/h2nnCkqOqACnbDRx34yEqdPsGe
vOrOh9SH+z4YbTpaoOgssXRUjeSgvHIxckfre9EuPrhAlXFqbj6BfoIViPKeP4NoC+IzP90NikIb
Kieuf77aRW+I+9PNFXFGihpHps+2R0Y3SB9M6I37MArMhUTyhl0Ik2goE8Fvo+KIKGfepFEpdmp0
3EIXBFTDxvd+BSm/Lx1ZV9FekuDVFS+wVU4hBArwRQ7ZM9A4fQogsS2YVhGzioF9R7wAA9cZisv0
o4xFVdBDey0M3tFtSf+lUYq0cVk334SS3ERx0cfUaJdraVeblRnaqDh+P054d82jMjlrC9wVb3WG
3kwuYHZhYWZl+YV5Y7EO5Vbekk8YcxSkzwq+Zq/2azVcDqftFOWUxRkn8EgnZbXQTIT9A/98H5y1
dYhBU/JRCWbZeJi+5rADRelr/b6mjICTegPHxsPyemVl0AheciKL0wME2LWLukD/lVFItOxwrAlg
2F7f2DvOua6JCx+gwGuMwamMTHIQvxgQX2yjISqCdwvUX2Jy63CJZCcCUeoVorBvtISiJLFb+X3A
oKN7gQtOggpV9ERcVbFRlTsLdC7YwLHu9lgzVy5LunZqfKh01EVW/mNlfSK6QsCdgJhC3z0sc5Va
GWxj6+1Y6pgrkxfBxIaeBKkRbkm0OfNkeVJZl6Yzc0Gj3X6QeHN4q2hFRj03g8iSzu88xO6HWY6l
HgePWXEG7rbv3F4HqsqGZsE81PaCMGQtxtKR54XH2ghQwdm7MY8/fUapiVAC1ZqTZ4Er4uBmU/uE
9fXOXFv5lUXEDsjLTs7Vuoou0YtgWA8TCJ1EWesAW+1etQJmAxbDHMFB8vjxiNYx4u/wZDBLOXBW
/HzKTbahmUlH7P0v5qMLTfCgrVO9h3elr4NAYjeDqaSNOgEyPfq2l1wUTTO3lzVKupqWqpX8e1+B
Q2Xetng4fo+Wh1NlDCkc3G6szj0NxiQnpIeJZs57XgjY5otUD389MWHbH3kP5XesYB34LbBGYaCk
AYi5eVOQunBak65OKXeSe91MADALpJxSO2JbIPGyz1BNl2b7/A5bKyFBRJFNebr2K0kTn7Z8paWP
UaTkY0OfvF6eSiHsBvss98loOTESaWu22b74IMAyuk5vJUn0nkl3dismzrWiofPoR0n8rM/jJGOm
ymEZKyWFKziVwpC4qHSAYP+VtwB/YTOddex8sQC41rlGWJ0SKlJSgLyzI0c2BNTV4zUzUskQ3wVy
4wBDZpe6Z+qR6Y++cX+6zx6Vw17ryyCJFRZrWun9bv8rQHtJQEvZBAQa6fBPUn4ek0aLIUin5F7b
KJnbdRQLPoJHvb32CEZO14Hi2DZ7aV7Q/Us55TFGHmVA/WpLox6sQ5XEArtL2Z7N6i8X6fDZ1SbJ
M29imXdWQwQR1wn3UDlJEJykOVvzBf8cD+Z6z0t4vsMTuUJY8f8YLLDmsg4wr0P87Z9lr/bmjivo
TNHQt7Ty9GgDYuGTLMOAev3ieavtB5Du5rEvZLRpegkYfHfy+eVSxYXzNdm97j42NobuGXoFdXJD
X7nQZW9k7MkacX2neZOAZ7iH29Q2nnmnWinLmWC2GtgeKnKzxhjStiCa38bikHYFsA2ETizUgzdb
aYlfEXvftCJmEszCHS2GThUjkKb2T7s5GGv3KRF/qNCp3Lt+eSln+2p1JzuRE7d8V+OBgd8KESVh
h00Qp8Uee2UN/AuppGWwH9rwtP/u8sEXn239mhbjsvPoRPB5venjnVmcDor5DDmWcVollPl1bFTc
3siFix//+9JMjF4bcur97dc3RAvSsf6bXOi2S/nJKONepiWUPT6H5UijS4tD370Vvx6cfObR5Tqf
yvQVKJX6Sc2HZD/9liq/9rarl4SVd2YzM/DtX94IV5/kHaSokLecQselEhQx6aNjHHS+7IXE8fTa
2yOublX5cEInupeno7CWfylmA3dflg74A0F4fthq9pNKOkpdHlaztBjMa32x1KEgRUOYFmUbSpRH
HE/j8cTBVH9c5RpqFCisLOQrWXY+SokQQ35hWEZnSjXhd8tBtcdh2hjxOEzXaqa/6/Ftea5ganoV
kayQTehDNhhcpq9UgCk1yknk6AoeTL5GciLnpe5p2c7F2aQLDdNHk6pKPM1/++Ow5/SDRDb+Vga4
5NISok/w2shDvxikDjXFw9p3epcu8P1v7ftvhSGmF0TmVz6xqyLGp5DwkKuOtTQ64BHoXCEyOPC+
rxQroD/sUIXvQdbY2Tl8sI1rAC8TP25cYs8gfEU3jDt7x49u1Btg93ElFrQz0LOo/WPUIkRUjWL3
nQ8JzHpNtmq3xWTVCiDDR+YuECilvsQ/s0wYwx0s1+zWHmjdapXEtGyIajt2WqdyXvB5wV5aSyqW
cbAfwURms8rdRPtxxv1Vec1/y7R3eqlr555NFbOkkEucxHbqMdM6X8S5uENFNc2yhK41f2+W3Kpp
flUD2wfnYI0jvX+jxshcSmLfAv8+QsQawUCjqSSBQtNinCxrqsBnlXIAtMl++cuXzCf0eykWhoP6
JSGRIqLdKqvn1KDF4fhbPtLXLpXRGg1rhFgdMyVNRIWMi5PnJUyxkvAuOSeql5TrJFYUZ5AgWtzS
YnQA4NKCo0zIaxQyMDimoECfFqS0xKtJmpKfK6jxu6pLLXOg5DrOv71J+agbDxjtCoS45Qkxqs6s
OD9waAoxYii0RFzh0p70Tzy7+IvrK5XLQlRE8hP8smzgPaDxVx77Rk7H85dvWUU7CDbD/SYA2gjk
iCGnIFQmuzaMKcXNVhrGXoyhMnbjnAm0bMyuyTxB29FhmJuj/aFEbJW/ZB1i/0FmwrwVqGKxgN7f
OMtevdRv+IeKL/6I2u2J/4tSxkocllPjff+IwHBXlzSRw1chpaTCFch5ECJw1mw6pOR/m0GTuh5p
pS5n1+Cl5A8PNz8Bbqo3WiGpMeZ1cL7syNoZRqvWLyOZ6R2LZOI2t4kctUrSR1FAbPUVzHov50iF
DF3OFCWOjXoTVmxcIcQ+r5NzuIDaS/QyFoX7oMIVLUTmofuwcIO+Nzkr2Vi6U/9bhBS9UqsmR7OO
Mpbr6R+kNujoSyU0oQi6qgJXLvtOpExe2Ol3rSYRJwuY30JZCxtVdIDU3swuajOjjllMYJ6no8OS
EUSKJa9SNn/NFRnUm6BzuxWpx1TsR9NoChfBQlyOeioBKccAow1CZkrd9Y5Bwy9Rg6sFs91VF6uV
y6YR//lSFj/FIjcNAVzloSh3g64AacCNtHNdsEP1xlbz1Ii9701O6wrtEAYI/7TWBDpxPSEeVo9a
coPfEUDgLyW5OnvI5NCULJsRCDXkFmtAAIlz2zq+CedcOag80coldMkldNXpEqmF8nvOPyXTIHDQ
1gTq1enT/kLz8jtxeTQ/UAFsljX+5yfb53v7nmUMezD8WP/IeN7+Cm75mQ0oOjClbOrSi/7jd+V/
SLRk8z/hpN7MkCUY0RP3w4oNVAx+viORuw5RGGVu/7j+pq9QbdFqdM9K5JyM5UAr/sQy7cA+UDYw
Q60G/X9ftJ+sgbkDwUd2ns3i62uC+lEJQb9tHZoCXfW2Cd0yfaumrTorUd44qWlIXSWPwZ7SVJLg
MWOnTtmGCNlGHe/D3erDJ9WYFLAKSrSRks/xr2+Jd6j+4+aQlS4Mb1pRKYvyO28LVOzZIUJY0lrC
aBS50eH3ZDoexj1EF0H0AaluG5DIgEbOHxt14TZQdrObb8JgpwYAWdT7TnSwcJw91dEPzBYOhI3M
3HluJz5Pe9tolWW9x8MR5dhY4MkeZTmoE5zkVnJGmbtRnvgzS+Tu4hn7TShTTqCAMjMlrc7UQzIy
LAZsxn6sbCNSnhGZFy5CsctnVK5tn17Cjv9FaOk/xAlQ+XoTUoq3rvo/DvFBlxvR5ngoX6tMkAfp
JE5fy2v78uoEFRSiBzdTNXi1ZDsH5QJG896vGzcQS9+bjGW8DMolAjXAmkkA8tg+Yrz42H3dkI83
iMxg9MveQBznNF4tZTeW2uQGkLgXrdyt/Rq9mbPunchnUchj0Bs6j3ILqK1XC9EPUB9nSk3Hq7d2
NdFw6Qi/NluWGo6o8/VmCqo0/APfVeXygWxyywqfLeVYPmfuuqq4YFNaRFqdFNztmO3qQKsMm20+
o9xYowtu8/URbyP7s4vz2hn+STGx8D4UUeYRWRVqaIgXuqdhEIGFDHQXVsZYW7z7258dGBxDjqIt
IPf+yIcpYmnTE2LCj7Fjw242lJtanRTXRfGxhnA7NZL+KVeinffbKZOJN8siQOqRDZF6Sb8qyXsK
z7BgvGvygbvdxbdYRCW/CG685i9tUj+znd3LPTVwORoBclmm2hm3bYitjrMt0Q09vNIyiaLvRmgr
WSPgtbTdpn6GAxY2e16KnP003fdA2PB8wx0CxDQBaD3ZvfoREhQez6HrOXlZbPr6focvyukdm6Kf
tGMUHbcmz2jwvYwrduxOya4QdKmkjyIiCZVj9JQKvms4ud3dJH3q3+cO2LaJyP+9nm169Cyr24ae
pxOs4BBUSy6OmUXyFYNT6lY7CxdiBSHCyHDdy0P6+swFMLd1elZK+zyoqO6Kp8QYcwAxMbXB1K4a
VAz5i+WmKtEqfa0Fx3KF+fyZdis1uT4H1V4Wj0D37IglEN1uc3mVA28xWCTwEBNJDI5mjtjw01Xy
kI+JCLRnrUKaPt7SizRFd+LgSr+ntmsXUSKqUOPzoYeSTnfTjrXPwtIiAVvFBdfG2a0qGVIOX9SC
/XbExoMVAuyqdJ3+HQ96VPB1BTTnvCUfY+7tor3Y0J1Ldf6Z1SwssO7aLcigHc5gaxX/JhEvb9sK
d4WmFQkAeRj7K409fzwkxk/6PdP1m57vLbsXvsWx6YyCsScrvYewCTfeRRFZyE62kBSSA88jfUko
5KKbnGt4pUS85sNGF9c4N0ZMC02lIqWyEbux/8npMkn2ezk8vftLw8AkfF2ynNUY0kBN7BsygI9H
XGi7u0vI3Kiso2Okz8BrnW+u5FaCsPfGUvyOjWZyL9XFkhRD8fNlHT4FJQ3s1z6yUbkKRuEeTLRF
MH2Ox+Sybf6LLX5Rkp22oiuy3bE6lREDsXXxpXgZBAGPPUgErb8ugcdNLo3IjtSJ2SXFbDqZSb9E
FKtE8WJ+lpeXA6xjqH7w3AEmhgPUOL1VnF9tJHYcXTZI5LhtKp2xlg5HdYzZSr/CkQe5vA7+a7C8
UugdlIbkIIqAnM1Gw5ENuCyTOIho17cq6TPUYEmcjjj/4g93K6V4/eTMK3xh1qcYh2lWFbWaaTGC
sRUSc4wKAKUgoC8NdlPX/F+lGwEAQFoczgRXcT3iXLiEsiFWIJjJZKGIYJe01fWgKrCAbH8s035V
HTS0TSYxIfvIsPqjAg/D3L6BK5XR6JFiA6CMwqLIS/wTyIckKz8SeZ1om3m+eQrFH8yApFVW1oNN
l7c7FrSsdQYBCXTTlzs3YlBZGj/Adpug/Rqm0mhJ9+AgtlxrJqePx0CGqmests1gBfup0AaJJeK6
uuUkOEpRIKibaw+9X895iMRJU/moVWoSRmrm4gmtG8Jsws4FJ8MlFTs8EvltBa5zpFMrSvpXzf1Q
ik4FH7Dd9E3DUK7/ulRdzj8CW4N+vLKVwxUYl79MG8kC7G69S4JCqiIKKNXJLavsMY6/S+NE/nLH
PE+pjn10K/6WkJlUN/l06XP7a9k4jrXoENgZkKIpERwXLcKILrfUh72jDel1rxrP+EURDIpfuRyE
P+i/GsFUIKqca+gHsS+oI38kYYcHlDndbicDUohww2CE2SMLHnzzfGuYZ+5yzwMk/ZlieE1xYxbz
8lc3TVuXFN/aiV+lCW26TGScZoF2oQ3FgXQy2B0mSbFvMOv+GXuaKZijgNoeOoDksFWRNW9xzNvN
3HKLJaP34mo75rZlCTJiHk/23POykBSbv8jEcKmC1zbEiaNTN9+63L47F6POpWuxAnUloky7Ls44
vwKlOyRj8qmEelpEG5VjfSRYz1zvaLYOQcuE00fM95eSjvmJDRVuhGMp6SdR+W7GHflvwVJwsIhW
xGnAcu65f0uo6nXWiyElBk5p5+rOa1rvMIWDUKEw6YfBmr5NaTsJhKa8Y4UuQBYtWL/RVxi3/aYz
BTOu4Niz6qSy0PYxOw66kKSeD8nFPS9y9Fcrg4uhK3VrNE9W0eGZm5MB+njmwUe6ySYvl4wvWSgS
j4dRCJeWESvY6MZ+4dCtJWdCfzmLu1TQJ0iogKEI647xebrgX3L1xm3Dp2OUlLNl67x//V9jaLQX
PDCRwUaN8SLJXnd2IYYasigqNV6U4OSsrZ6Em4YoXF2TK37517CCL4XadOGQ9eJ6p7inWkCPYf3R
KNjQgtHZZXaZGkq9I3O2EWWxP00YobCkkeFMSLYCbk9BvP0t4Z+fetQ+h+MJV6WeDUANK99W3ajz
HeuwaxYY6I6SplUmAdu8imKqVc1zZSs4LXZNO2A2w7VbCjKcRmW5UC0msF7Rn9eDI32SbvmcV7yD
U5Ws+CHpVhducoWBKow4vBEJq0+EdNl6dHy+JllkU+tx5MapQsJ9UrTGh9yNJrS1gv/PgNICh7aX
jQVJ7PZuvp4SzZ78SIpjrsvkUgbE1EcOgJSmDiRJ7x4cpvGwffkKsG6iB9LGJQPs6kL0ZKC8KcSB
l9WX0HsivQpiJJNGoS7Smfr6nnggFrDhZG08EJ2r/8OkDLMo6Tnsgf3jOtiahN6jSsKJwqDdrLx4
2mGsSDBJNhDo269X0/O8P5BgaiVzjImm93SOrJRpK2Pel5c7e3W4L1hFeAacE9W6sOeQFqRUm+6U
R9F7RuweFyIavlulr0Q29cgN4T++WiXM3JsPaI+lB2jrXyNJDgDrkOjGI9EPra8+215tzJuEmr1V
BLyVnhBCPNS93xF9Rp60pGHVPDbsBFjebkHuXjwSiMf6n7zJPlFMkYmwx3pYVzSK8pTLELme043E
3kpa0bwQGq8Imckgmis8BI+2Sy1hOP8XP6MTvz8uX9ZsmZxdjDC6KSprDIyzAoRGipH/NYYqRam/
jCjyqxYB6Onrxw7SfOEJuPu1t+l9ErfzRY4JtiXtBmRXq/G8ms6vRySizeT6DYz6rXE+G28mbNfN
1L7JXwNIqcEYzHGSz+tjV4+iDXnjypIUV0PJV3CHLsu50nJkS9rp3X0j0YWANmUQhYEjZVlGYVD9
2qEeYPHb8fAgG8hvy53VEAkjfjMDtAEcdb0UfUJCD6EF5eccqFVBnJWlkyGXmq96dgUfJk9FreLS
+JbGTOq19p0qm2TOSO0XXYPEXpKbPlO8gi01TgZMF85lL6EIvk5Bo5NQ3NjRNXXPOfSyBJJDeSnb
9+gPUNJO2qfuvBh1O8xkiwK/+ZkeHdzbp/ATSbxsqViEn6WRh1FSCeuyeFLp5ZA2hkBZfGNLWYQR
oAgP04QYzFpjp9vGPmreVHm/BGAHn0t7E70cuhZkLpZLWqGyenk5LkFYQ+kiKmith7JNGnHMQiL3
Ep4EWtwdSdnML7rVXfOxU+rYnL6UbuR9jCgC9jN2ZvIaZi3Fu6U1WEhQkx1QKJ368zrGLW6uSdW7
RPvZ7sRRQUFKWkRC0U15gmk+lhLvUpZ+zxG6no30F2YL4on+ioNJd3I1D17sykwJYIL1Pnd5di12
CClP4l2cmWVj0m5/B8vUDNpz31QahrS0yPbPUd2YjdmkckSmlV/A78OS8AVADXxZTFG8RIWjYu2d
Waf2f7OPrCtCOJmzwFwRMLymDqEdCBKndjykA7zSCGaPuYIMvkZFPAQofqbyYTretoJqwDFm9dZN
jjHa2Y4J+1Aq9NvD3ewmUPoa8F3kVAOiwlTkF/AZAuCBPwwT8Ix2zO9ZvTQAuWL+MmPesCFQIxuT
dxVuwxVPJastotAr2LpMbH/AzHdaLar1QvgKaNuLS0fGHIFzqbsgPDNolHiBxx3xpigPA00IVB6X
+XsNgPr8xDaT4fDtoOAuSZbtU0UZicj7mpsIJdQ2xROfDtt+zQytpRbIvFUQGd3yPxcMIx4et1vh
bPsOzhftJ7TVJEo6Z2vEUv4oxvmZpugYPxKDnUUSSRz0AM8gyQ5yF7/O8KzzvP7HaFRu11wyBcmz
PnS4Flo5tWy0H+nA05qAxagcJ1dvxhL6ZXvNqy01ZOTIiGFUwClCuTFUa3VzSqYiOKfn6244EU90
9w4jKNallbHVPcZwAkBW6dKdHBSa+K/WB8cYfEnXcir8o3SMU/ZQ2XroonAPueI0iKoN3Mn288hE
g8tOKOGkopU1vByLS2VQS3eljxBRIIeSf2BVpbXrt8D7XUtTj21f1snwm8ElW8QWfSqYmX8tNpEE
EZi9PXZaJIbtbgnCD0RTjGYr3hmAqI6saf88qNgNP8GRPCeu6LIVZMX9HCuIhzB6F2llUu5MZvn9
5rizfxO1TgOsowoIkuT3HV++c3DsB4G7LsUTbI7H/tfXyOiMIxaYVdXrnHebT4gqh3O4nkknpQ52
96KKxWZTqLPAtv+sSFIM8TjThNjJ5XmCl3QQBJvbvNpNAk0XE5eVPfeYe2lXwD8Krkx7WlIUHw6N
6BQTYyWX6NkSwyZuAinjQMCG3WbVQ0Kzh5HKnacQHkHRQ7PNPYf4B0tdkfRxv3G6j7pk4i4JmrIN
G6QohBFk6NIOvGvUtHfoOFbCGuizEgzExD0X00jQPHG14znEKRPa+lQu0oMm+8IDfTIVEU0BF7eW
84kuuYkrRV7188fev6/jtwUySHuGfnmgp7MC7v4LYrXTMO/jCgtihi9OWZ0ZM0+WaKsy2fTq/6U1
c0CQvywod2vw7UBkyDfNL3QytFOLH8uTFMm2+nCPGbW7P2+gYz1GTo5fsmPKqDdvhQcBVSI7KJIv
OaTfcQjHhTYtayMKytTJIHQO6e7D7HIHPDbXSs9WiXUgb5XVPEAbl6q1XwPGOgH3T7s7fdiTSo2E
u/0UWz/w9mSC5lsUGMSSiKor2FkIOvyfRG7rXyHkkJtVi2gXhbwvq6kzJPlbdOR0L6t7pcZHPViK
Uv91AphOBXgGO1femEO4DDt1oKQEVH54pT25PVedm5brkwIk7igqKQniW52kixWzd2oi29KpJ1Mp
WNLfQwCTxxEnvJXTgqH3s1j+zlwkiT4fGhAEEcKHX8Ik6Zj2yOn2JSbmIK/04e8UmS+6k2ux+19b
HPG96vZSOCONMnX1dmkaOc+ZD7s9O3j5A0o0EMJxD8GI8wimNBUaTSwcG8pRPANDDuCSmrtXY+PQ
xSLKROCEla2LxMaltsEeKCYcGb3DXi2nBuGc8iTJaOT0RdSW85Gxkek2v8FxLTUSFKhiZ9BU6ybX
PDHa/hu71M07vx2yGXdbnEr2wFMxZuzIceUOuSW1AR7BHeT0s+wM1YwUojtJvRdSQiFN/B8Ziwt4
Og8jgUmnPkBSmsyLZiukFZo3uOkR+aVA8fooSoeEVBZ8BQxYRnJQOETvuYSWJzJAdCy6KVDbE1SN
j/B5hlV7rzxLgfNfPCwm+Zc9O7+/YsNl8j+nvo9i9z7YJYtnQytxA+9z0mzv+ydJhD0XejWBubLV
Bqt8hpmSGytvMiuPHTbjy9NBEFWfzNPhGEnJsBv8VbDf6AEioIlQV0dPPOLrXiMKmHr53Q2KLa96
tUNQtJJMPHjKLmrb2aYs/yhstW/npiO33BviwKAXpJoelRn+R6gujWsL/MigTGuMlhsCq5vTsxTh
8O+ieMJN1r7jP7CrzM8YpLgmQoFc4xaH5nOXdtMiIoplx3Dp0C9I90ajO+toDKC3jeA/LrzzV3HH
r98FlaDrKLNSxPzhPsmNXNGTPdWmr1I58IdfQMsW11U5UaKsYi7E8LRrr497kOIuyzHPIng2Bz3o
F/KS+lR10Dj4wkdyIExWxd0932pPB33X8tdyV2iyvChoRaLs/WpmchBNG7d35gxPDthrAMHywFos
e3jv1cKzLPM81t89oCOMU4+vrDAy/DaK4GKGa5eDj6IepFQqNGPRNBBJ4WdcI+zhu/F1PfCOBOTn
aOZ1a5xMpCVgrRyqb4C5U5mF2zkQGrxVU7IhAZm1XHeAdm/GgoND/9Slpe1riE1t5nbrMdBv85F3
UbifDEcE1yKW+yzw6rsz1TuHNGv1ICy1sIfJZYZYVMO8oBUuO8LwCy2X6h6KofeNj+BxtqlcXxOV
3YsZdV5ObDswPpfdTB+pM/+d/Ti7TM0KV1jyE6wvUwizb4ecg82VsOQlnLwzZfhZyqEH5Zex05Or
hLWBnhQcekhb9b8AV0uA2PnwBXE71lDESdqFDTHnmCrrrnG8GkEmVQU4r9+EFQuofZaxJZdMwa73
6pAMPTd+KwR4zEWt/DqgJ9Pm2ycbwHUYSvmAF/hYbJ3g7Dntb5I4i6QWrGWHRy1ySw1I/yTkyHuQ
Wg3fv3rE3s3jaLrTwAG/hyHnh9dZX98/MlwbWNcP7CnQBUp0NDSLHxt11LyO1L+nftHqoJ8Oi5lR
8IcXWgFW198a/M5UbwBCq+hQQthg8BeMMNQZ2BvM38KBy/eJpUF6obLpu/Ygju45VL7s8bOPJcOw
lO6d7bki/dTvBx0Xn9+HJ2WE1lY1daAecQT7eSffoO/hKktCcAw9dBxA0E4O7TJloU8o+JnbESOD
jPKJcbn6QxZd2N60pERyNGI+vEFkR9XrDVJ3xtJfPv94+CllOwuINPUrNHWA2nnVr7IbIYWiOtti
PfxYHD1PKOswdAG0L1+/DL6nG45PCdR0i3hHCMdNH4xehB2qsw6T1p7C75Zl/t4+cWQymBnLDbar
IoHf0JW4hmxWYrCCiopb5gs+yTYnWlFOqRvOh7Fd/zGJyXQL5NLq607LB330597lao+NXX5covoP
hh2OIb5UzhISeJ7KSptNoH28gLCmilBSUVJs4EiEZ2HfT90iTRdWIjXuff1gGelD22A6cUDR/Zqr
QWlI0AbpfTm1H1nKn/rmh2kCtiVvOET2vLEYqYiRhQjMstdbNSW6mA56muCGIKqGABs35g5Z4Wbc
IjncLPKf3JjNhoCUqtO2+n5JUPVP7ziTiuAlucCVR6Ounh7PpxkaorcYpb2W2eipn0wKCAt5rNzh
tR2UQCQdnMwLRuFHA+q6+nzkBQCBd9HetL9VbxS7y0xWUYcD8NAMol8kS6NDxApGNHWqkAEF0T1m
qwVz/uuqR6U8fw4JorFLUf8ynnKkmeohqETI0FmEX+SV2B8IfA1x4dm3GKPsCqQONAlLVdJ+vABn
SMn+cQ5nbzbClzKSxGZPQDUsN2L4evBOuhezEeDl3TvdNTmo3ih03zMxbU1emBojZWZXbUAs7m19
M8NkPIo8xaQbg6pRELH6nVRepXtCJ+BvnhWvkV5MfLGiVatXpxJlXsY5NVCaiNR0B2xHjGis/FUf
cNPzCAf/vsV0Pq2GIxoa+TmCb/EAyjio7W9C3sn8NaWGss78JWXH4opVRbAkYC9f3P0GKlHgEGXd
uOTg5qCY0T8QkM85WFMCHfxMzytt4YIl0I2rFZCzA12OoN+mDcpUYkVbEW7VrfI/2wxCB9uQ6XUC
nQKVZmkpSfFw+I7ay2xCM5x2wfDqoUQqMP0WlA80I5Z+2fFCRKqNyQ3wUJv+yC4C+OoXzM/a4F+B
6ep1y7IzWSlviZa4no2wxgF2rso/Kv+mJykLpuaK0eJRoSv7TKj9Y82qflS5CNWhSnqTQJKS2BHa
c64UJiG30EtgnLLNWt5bgDcQYk3YMToqb5dxut5wga7qUpInzh6NTdOOtJvrRxcyItJPlpCWTMat
up2zd52hl0+Xy5Bygb6Kda5nCX8JwZZC4HjVXteM6mzIBlXDhMx5pl0O52iz/c/nPmbWeQDn/yyw
BpJZvVD3PSVb6YcGDaaprpcR0qIkjSwQxE6GNiDiXUXiOUGnFzbhD/fj2CTIR0jhPLVstuKL4HUt
Nckw6NPReJFw1WQiPbLLJ1JzL+roLtl/m33QbhjC5qaxoB9P2uNaVafZHspoT+3FLDyvLI7hBals
m7eFn8yiDSjGl0pxXFyOI6hRMtDr4KLQOZTlAUpKRDAl7hW+EQSIgHMS2RyYjlS+CI+cZZf8dbOu
oCsjfoHfIK2HAu9uqyJPZEe+MziybS4NGYjSvk2E8F0CO39XgakTYpvBuZy8Zieo2nanVL3BdypR
8SeXkkDmOHmp2Hx7bOuTLGDTUVX4fuUUK+ooO3bDy2tgBCi3BS66eIZVTGHctv01Vwa2bec1y2ed
pSG1hQuOen6KAzByhW8//NTWPcrSKL50g7cE+v9ipLlpeOC0KoFI1PAawQhGcsbr6WN7oS2mNplq
HFKrpNve3KmaZt8/h6v5D3n/Ld78nzrENYXm0FUr+b1ziskXZtu0G39qLoBqTu4ds5wcJzZJuBB4
Wkdf4eISXwYdxcx5tjL/5FKmhhnkiKJ6hKsfmVNXxY9wPqIya+ySb+KLSFVrbdTcgvH9T2W4Xji8
2zbk0g30huVPfxMfltxdwRDzOKcSHrzsGF8KpS/Bgjbr5f4vS5jYnd1eLae1hmrzjGkTuEpf0LID
6hxqmFXvLcSQrar/APWTdnO+zyDhWl/XOHoLtvT34Hqa1H6rR3pNqFJHS/wafWnwG4oB1SzaKngN
IvYnGWjz9WchcMyLIW7779aCoAiDOlYRHn8UZz5+8ZYn7YHv6QSVsDqVKQJAx6vyTKmAPtjStIws
EaO/OiYeRxBbEcuxYbBd2gn5/8CulGuCzrTLU6Z6z9YFyu9mTcPS/tuceXTdb2Q2JfsT9nU5/w+N
9E7A8pfKXSITOmwY0xr6GYOI2dW26dd1RlYcoQiylO57YV3iwfgR5D3enGbFiwUAkmp59Bs3bHfq
oo48M/o816tsUy17iGjIWiV+j734GwTTU/JDrICR72uU3mdIcjiHZhwspztTvfNRlyUWxUyOR/Dp
o+hCJKtiQyolqnVqKBT5j2tU6SdUNnegC4qGyOOTsUU8F+pqT8Re9R+ht6TNjHRMjd21AQt9XbYw
KEYAs2d8uvN6ju33jh9Z9YSQR536wV8RvSdptw+h4s6Sk1czWeK0eLi6hhRWuDTDjR6m43XZT984
2a9C+h1gmARTkQzPm+wLoRMRfpgHBbbcOqpNT+P5teV7czAuEFLSfIKSxwmRqqudHePBruZQ5O1T
AX4JYvm1g7FXSAwb7EXu0oa+7eYpgWcV4QnEx+Nl8GfKAu3jw55mPUFedsrBrhEOTBFx/863VXjY
omebsfwDhiLEZtz4O28iWBxx4zKbsRFvQdttTeonaof0hCyIVxvU4i/olHfY86F6TAgB21vIRAyQ
1d7WH1axySrzKMwEY6fGyA4FWfQLhZ6nAeG6qmmhjUqvsBueB53n845wyWRzqGpeVUFEtFtQxq0Z
IfYZBwnYBBHquCHaOWATCnv88K3V3/75Z+sYy1qvAPKBOUhtZT9XzqGyBcp0lIPNpqf+xp0iPB2J
b1K3D8N+wC56qjdbou4bD4uw77V9+6GOgac6/LMWCKRd4ZNoMIgK7j4O0pPjp5+ItuXVfHeQ9fOb
DFuVF9k0WE4dp744t+cVLSdv5HiVCHBolYk/8Q1dq+wVV+L5+KxKyHyQgR9te0SMtD5yDI6qWF3/
AJVizZw4izeoTGnBvptIofcF/Gr/bzwnVhTM6c9UfCbmN4e7cV93jqIUip2mPJLwMwMsZFZyDLCB
uszTXs+jJSbCZ1BF9qPUwTe28uwarsd/mek7PJnRGmeWBQwqa39sc3FhZgyPGTkntwSS7f+985U/
NkL2jIIlwPSrHpr5NV6+8dI3tu7jdGH1J0vbCbeWprb2SmMWOwoaqHalYShypuDruFAXKgJXJsav
DJhPjYnjVlaiVs/ezj0rVxDOHpHn2oryRsQRD7CEMtigY6laaavjj9J3WFeRaGc12gnjgRY9U0g0
Glih5XL0TJFZHtCJfplQ5WBjLu6keDdjie0iG3lfpiqb30rYL0JtoBScEUdz4p74DH7rjpFpMu5l
2FuQjY5XNBqwWC/wfq7Fso3oXbjji1ud97TztnolT5bHYbZ5u0o4PViqDg84q+3L4yB1MrR59WRx
NWkI67b014VZS7xLfhLIs1GtRtVzeqk7d7/putV8ktTh8T6I5WrbwGNWQKKlvsM2o5BCpuvuA06o
tFfVKkWRF/jggn+qIb7KV3hiqPPWXxJhuPQMBaUN1jzPLdzQ8gdGK0MGMSdG5dfKGhQGl87xio+E
0ixhOIUdtTwPUKnel1S8HNeNtlmy1x9ootj+D2PRmZER+m/mZGIph/NCuyrJpH+FYGFzrytl4VdP
tb1kZu7ctjOoddOlr0Fy6KSq52B7kUKSMGrqrxNkhhH6DOxzpl6pWnZd5B+NqE+N1e+/uJ4LjvH9
zCJ70kwAGuZQ9qgOne1ctUHt7fVDzptIUuzETC4EldhAS/8x9x8XawDJInAjW3Q8VxPBzc+7qj/R
33BDur322gcYA6hp1vqjUvuU+DLNKk13poX78LZ1l4UcwbUDXM24w2UjoOqUBRWLWb/+gJqSMlav
Zlrick28GuGjPSqzyVJ8fKSYXHJTCLCc9Zn8TTZ6Mms4/E0T2ZdTDhSaSXHIZMDzXC59HOt1fzGf
yy9Z7QFIeWgRUjl+yhRxVw0qM6GSFPtRqXZ+3p12hc778HTfusPcqaIIf8NJSe1kgWyfdZnBnc7h
8ph9I0rvPSSvRNiEiWTK1+lO4cYXAPm0fAdcrZNzSQlXrOAxCETYWtNW1qGD7eC63MHAzdF2s0cR
PiT3jbHdThEeRke/rcN9QJm0cVcqLLLUX9VM1D1bd9NmI04rVZfczue6K6W+anqfj8PNBo7PJLTW
Ocj7a188G61kAE0fIn4o0+Q4SCDNkzrFWsgTvYxFMwwWImb1UhuUdQqVH7BJp5XX5JgKmZjhR1Kl
uIh9jNIoCh+sITWcZDEBpeECqx/N5k8p/AP5mhC3PBMNlvRZSKKVQlksljSxgvju4MyzqDL4cLDc
kKPPU3Xwu7DSD/as1X8/oU36mMBornaKrpa6ZnL+kPP8NLXpVi7bIiQ/eHoKXi+7BzcDZ0XkDq1a
rRnYvwwJlWJd/aj2VMk9bDLeuHBXMcUwwgYjYlEsHirEhLl5k/YlmHBhkOpW8MnKzcj4ING/Jou3
I99m61GFvig2FRnPRl1WWoosdh70/boWeIlz0N7jyCnkC9xUsLZiEnX/koB/Js54hjCNW3dCilk6
OrALY+5fjV/cE2az4GmWdodTG/hSNdFeJWJydVR/gDvly2DsIozeXIo6GLvltjo1R4MGHUjKw36R
FICmjadndWvWXig++BRmXDrka9av5CSB3HD9I2m/70nCCjib5LE+bjWFRhmhWSLweXBFPgQXzrSV
I6TDJZJrDo5OiUTEBhKACotkW+XbDOQ8/SVrphTpLagnueEdrYGyyOg15WUoa5XqrwiJSt/fIJ9R
ahdete6O9CLc0hPMZVntCjJ61eO/qYi/aCYad/1Ze8D4DGtAaRE0JL7IC5sAL7h6NmTKpCqAA4f4
yPCV7f3pWN4ZOq1onBDD42y+JlrquJpdkUGXs4kHmy4mU4X4r4cz0LNfR5HcdCqW8CR1uAAzeOjU
CgDn/Gj9WNcIFseX+sAmxbRBECaIPibP8PcJ6GSD1RWdatgcCHiUtaXAtxUZSe3RqRCymZgTMiRg
vb6QK/74+w4vvGX68JPBnyyqpwoen1lNg3uRynDCegLLYiz/CR/G17PoqJfqTvwNMcA4PO3dJrmI
wPx8ozUKMhdhp4TOnboSr2YR3cAgvbUr8wbitA5vU5L1fN1H4mFCi6MIJEFfr8r+uuYUUsFxAVxr
L5ziDajE7n4WPRUr9sjPV0R9/ywuy5/I6CWffKcQrN7PNepVY8jZOb6zzX9ivnRx3A1znJvLewV/
4BHsnm3ioPF/7I+dSIfE9XzFJlXB3BmcZ/80mDMfNsC1YbOHUum56s1ENLnAaomZD75zZXJ7rcpX
nA/3LINN7RH8hr3nPM4/tGQmo6mom75pKAOJMVVR3J9LUV75CJ25KeW1R/suUegVqf5Ne5RIFH57
pyrY9MoTvyb3RzWk9Z7Sk3X0DWyNH5UDKrxysoqDglQOgiEg7OYYHnAgIzRKY52TBQSNfpYcEyqP
nwi/khHEct5jFQijccTo3r3Eg5vGok/WGb5oR39imvTR4i4IipPu8nlvj75rUErlG9eUXnYt9Hrd
Q+0kfDehGXEgPThwrlXwskm1CbMHeLYqiXyxtWz/Rudl+BxEDRDYfMiZEAnt8DPBzT3JScQL/LJY
j39UbwPbIjkBASXKLZ1Q6xkOTaz6kE7Bp2p2Rg6Tr9J3ek1D+7cOYc6cyjHj2Wx8k4kEq15Q9Sxc
eO19zrZUuS3u6jDzNvNalFuvCD/hEUBRdv3RRvuC5YWepVPbPII3T4FWQYPBI3B8bhkBdj9mdCne
DPVG5cjj4ikCLhDEQy/dgMbbCSEVWuP+JXijhEbh4qhPHvCql39pGM0y9IGCn9qIr73ld+NQzR0g
6dCEfwQBtRxnN3Q/z4s640IgHS9AVKQ8NRedDPOeSbknnW/9FcHAlwaAXtpCptCH4tuIO1f9nNFU
eijJMliPH2fZcWU+Ieq6RGWldkkpaGu+gqzXm7uSfP+pV/yOv52ard5+Ym2YPf53zPVakSlxc1HC
lWxXGFDacsVFfxbDJg1Ugfg2LBWSlJYc82P3ehPywyrpfUjyXtJiPHUr9G8t7IsWJ1LXtuuaj9km
/3ELxvwf7UVi8le2al/6zY9Mxt/fCr+kGRNMD8fWI18euiRr2sHs8ste27U1gTUprQ2J8o/3Pood
pyhpPzWZhhQ6e8Jw/SaKmJaUMWOSRCqAdGmxGx+lR39lEHfRZRsW0NaAc3qcpyuQrVfnEUWw04Kh
NXRfcYrVvhKBs9wJGFUY2PQPLJtxSrY5QUGDRDdvNuDPfNvX03Z9mQEpm4K692ZAEvZ3KgvGZXiN
i5kpbAnUdOkNTMQYKSCdNVCkTTOW6VjeSiPB4GBvuCCGjAlsQvLecPhC+o3TdDFwAcVE6AJIWvGS
5Yeag5R9ZPO6WXB2n4e8Z1Zb7QRyI2uR3k37lSEVa2GsWBQ/rXNWyjCY72jIJ6rAvtiL6ROy5RN/
SHqGRlgTLtC0S1M2+d+KbwmlkPmdh453IfzTk6HS/Bxah+c3L45fOu7jBdUkDLDcfOtUO2HRMtJv
L6SlchxedH61qW0ue58W8i6r4GvCG5q9Ck1dyRZpgBna3tvBvovKq4MyhU40hYgmUbjqH+f3nNhL
mu2LbjiMEuHCyOvYhvCG4t4icY9X4sAMhr8r0FBrOK3yE+MHSccpXokyUEnNb4TztCwB4c7IRWh0
QQlbnWm1nQQYRCkc4Lmppco2u7n5B2uM9RPFRZgY2cfmEJcVcuzabDXht6b8vWRTfy8EOSAi+Lm2
P4z0QkRa+6LySAQ9NnzrXy87G5606mDPhmb9iRF6LZ+PeJIrjnFQxPUEjA4C4/q+4qmSpmvhT8qs
AmPODPkw3iqeWyZy5aGDTvbdRrKc+epDvByVMJXT4fJ2pQ+FepMs9TfutcdduMDPmdn1vf/jag+g
J0AG/mMK3zukzBVoS/fa+uU0rY9+k30HF+0H9vwckOauVLGM6ijFRFAw/32P17bOTvAUBKK9PVQi
Lu2JL/Tf9Kq/Ut5C6mIY5UFKQO/vO9R8gzawYLwl9Ttm5gHCYpd/i+orLqgWKiOxZ4VGQ+sBtcaq
IUJnWfnOpdM8pI0YnbpsjdGMVaJCmCxAXhXw9hBRey9wiUrlG5HTdfTlzOLjmgVBS5EJfOP4gRV/
0T4DcsdiHlCmMjmJO7A6qDCK436J05SFhwCx58r5qeWAsRDN0GR/ralWLl1NjcHTPa4zEJkmH9HX
2JfHYWSkIwbmb62+klUX4k+23cl0nZGn8zoNtmlo3nAEe7yn53+T5EdUauiQZV/ob50ShpRYXRiZ
2Bx+BlLGATLLpaWabMep+nBZo6DfktRNKNcLFupzyNaMWBjGBfk8plLmY14JmYasp4lP5H41BAPV
7wblfPjSBwAG284ghRoTHxUXaL6Z434q0Fdlpq4MSOnPUKs/A5eq3wRV+Qq9RzOT3K0vnNAu4UMo
qCs7JxIGCP82rG5jD0X1aFCxqQbJ/WFpcYAT85LaO6CwmhLPfScEim1fvA37d9k3vY4wacaTpkLz
otFmpF04eHfNwBE5Isl6DJjlPRY/PWP6dI3psHqpwNCdmibXL8TfB9bwb10oqPoMYL9MEB90M9nj
q7HdMyh+6TurTJSpOgoYzhgfMnC/FugaNM9pPkaXyKU5Dih+R/ROSJ285xcbNPOp1rYq2hsH2PRT
sDwpFlyFRHapcOUHvp5xZk6+2jT/l3IfwQUvAPZcelOR+9Xa/myEtjFt2sEDUz+co3I91E1cUL9w
e+pfVzuX5lw+DQL5LQe13g/uMctFRAySakWyTH/ToYdDxFmqJZTk8Akuh8oOlij/hiGzPc0pYBPq
N5ZOXRBgsP2bL/QOsAD7ewbs5Z/ipB6S0Q+duct22yCMmUwyaMNhQSobFt4I1+9VnSJrvSAqtM/C
srt59XdAPFFoCTStK3ETJdCpaiJrZWvsoYAP/1QrTDO+sFL4s0ebU7q2ZjbYRWiBHfvKS1HI+u7m
1tUQ7naWIc4MYYHJ9NzD66ef2uE1oOi24uu/2kkw96fJmw0T+InLwTQRjErqfljKjTyDXuo78yi+
eMM0LWkASzRx3w7ldtTyvHtEra2D+/4i7OGXoNMbSFtyAKLEUem6VcB8KlvIAzSWJLS9+w/ALb+6
Pa07mfBsYUuzpJtzjFp/2zAJ6WHzHnoapC1WlaMBY1dBLe8TgKsE+vgyCZfjPYAL8gL0H6E40bBT
TG+dmD8J+OS1bzZlgZWjtqFtT9l8k2ujun3lzP1UPp3xQrg/JEXpr/5CTqCEq3xzyaqfBsGqxt9h
zXL7t5A3mySbIJLBzNs4k2nPTeBmNW+536Zs3cEhYXsu0/ztW2BTjUL9KbiDhxj3KjvH7olpdoVA
QE4CZkaMP4ANXEz/K8MTuZ5XeopPLbD6MH1tc5p+Ghpwc8Z55e1/8/lUkEvkCBVr2yRpPOw0KR5g
DRLB2tbmBcjpUtjvE0jxWRY05ObSgmvYD44IzaO4xZrqTYnIFr8x1HKa2yuLaZWWC5kNXk5vUmTz
dVIFc1fDJvolGkk9NeCZAjOyJj6y0qQR0YA+B5ZDIXTD6LS0dH9gWMD0ozwIo5CDOiC2S9PyntM9
OP11+twoZi0D4HFvEeACco1KZ1Cu+sv6jAQSvFcjmNC9FpwhzR2ruMTCrD66uD8IBOmZBFsVkv64
yZ3HbqUs8kCTdQmxq8mGwyTV4arnxTqEKzJunfaVMIc/3g5yO7yC4Alvq9tB4KfbjYayitH2H26U
gDR7wa/vmbZIzO96mjaDRK7IXzSW0l8IXbzNaMcl+MXP9HoSknU5cdzg7pXFTKJWuC3xPGzzjkc4
1tJ0/q/MqHW64sp/MWiUfLe3mh8ktQKmafP1CGMo7Vly1qlIq2GHyiodPiVDs5/J3CLXtrXVjsZn
XR70LueApj6DC87eR18hYQwt53w1d5BIZoIbhNrSu7WnUBFlIzQBhwp323Z211Xz2/5+/DP8q/43
3u5+C/gBYovD9uGD0t1Gtv0QDCL9bLaKsM6yYT3MWLloeRxd3ADZPOKop7LF04YpsOWqp4sfnBwE
hVi7GVb4ARSMy/ODh9rnI1YyW4ZCVElub6MyKGkLTCG4JcuwD80+q3LVjPC/XAC+bAvzElsBWaT3
MDVSmkIfHWupkPyQ9ZfBMP83pPdQU9S2w39R1ZC01WNRl9yWTVKSEOqFX5CgYf1jNJPW2cTPxmYi
L+Dzjoo2+0l9fe0dw1Rzb3SoHq16b/xW9+cP9iB7u1KNE3o12kR5BkORo9sJ2T1qcFTUs1M94kON
30+KuW2Bg80sPMxX69mL147E8HgZ2kS2c+Loc2HHSVx/GAYWmutV9TNZwfa4YTjvDOWTqWbv00cI
6sz6iuN7Xx89JGGy3bwyYiN6szps5YO9VY427nOCyDdLs5GFdGJIKImxSq7fFVBUTyCheQMfYrfD
1tqSOk2TfqopX5dKg7pvdG1gjdNrs+vcY6MuMFxi7rH0SDWLRGJchYEPhLnaeJskp2TIDQERJJBS
yEdL7W7/KeSSaFV7dSYMqpNw7PrXlCtkDmoaHnav+uuLUi/EZmL21wrkNf430SCuHUbqyzszNQw3
mV483Ke5tDei9nIAfzGeNhhVfRT2wsAIwT7iXEIncLa/IaR+/ZhALZne2DScCCLm62NFk3GHMvD2
XWxrRRLlGVZOKKXEoq1t/3KO2kxTTVROPjmUlT43PnbihXne5S23MuPt3c9a3kPPIu2kZXu38BdA
LrraMJ0ZqC8gindIDnEY9kMiV1JhKZiAQoyp+oG/uWnK01/fSZWLVUhLFSTcYNnx9hFWL0sIcqPq
DNYZ0ohPcmakHr/twBA9eGAsdYfG8a9kD75CFCJzTDqedynmIcAT43daor+9Hn7d1KlnYmDniy3h
YqoA+EUvAZKnNre/Odo0q2eHRlbuYxlXd26z8MBtB7938cD/HHTF/t8rafxhVUBuJ9ZlrLzecJ7A
Jw/RWfrAeKhAQtqQLoWuoLInJL47PrHCN2JjwBPokkoYLRneg1u2eQrkXxg764mht4MnijlPjwyl
nXXQ7lkmRh0VqPseL1z62JPUBQzWTLAql2IGIWgud+ptK3G9vGaWNCdluD9qquLEGu9SibxOcGPu
xiogWVL/C+FdZ5xFYL7wjBPlpTMHIix7t8q2411Z2xWd2lgrLMP1J1BMrV19kaGTLSc8S9Ylu82Q
wd06jUEPBCceaWQMcIOAoLpVfyKK2m73rvE8UpC1vV+XoqOj//TZrjqSUurOVcCd+QepO8YOVF4W
6ibxy/FwfUs+e0AJ8lnCwCoym6m42nvh7CDjV+81D42ggy4XtB5f8bxzfC18j5o+S1W9C9n/HQYF
5IHcjwdlkzqgZGsx4KmjbohboxmWvjm46PVm3sZbq/gOcM+lFAAFnBOV2L5xHMAZ88P2hkpamFQH
7MqItIROs5iacS4bMzqZJTsw/zwhIBspET0ofGXoyvTxutgH18BFTtR7KSV63ccyJkWsKH44dj0T
pZN/zWs7bgPJIh3U9W0inCVsQYqOggyGRveLrVZEtPKC2UuslJda6yzKfoEdRTInmvjxkIDwOUFG
SWeL6+JoXOTnQZ5a28T5eO15n7K2xOdHiYoQJkZUV32OvJA29OlXffBlexR8/8+waDQQqgyh3xn8
8WFQ8AB92HouUHYxganN0BdH10r7WreEHGarvi63XgbzKjgI198rjRRM9+LFl4dFFdl5CXtz4l4U
+5/kDQ6Vt9Ty35fjMiCnmR/MjMXDDXHLMKK2wvsuN1/nxZFulu5CV4gbMuf0i170zMKxI7v6VKWR
Fi0yLoA/zy/yeK/Jp4vSI0fkGdxPN5bSsXDHL8dwxkAHIZ+a6gCuwXx4S6DiPPf8ZZnLnxxxSIop
CIivaCYQ7Rhe51DT+Hsg+ioj/3g/lVoZodjE+D2zT/0NNFJbbQhwcddVyh9ZqKT4F6wA/vtwPtmK
DLd8vztWIDFOIawE94xySNUEu9TNkKgTy87Pvu7w8RsnyZbMngxgaDh8Gw9Bwlf2NCD6CIWI49F2
cQ6K8YaCelBKxwSJBui95AnkpVG9/iHdL5+DXUpT7PhEHbsA7gzcWMO6taodPW2Mmfx0Z7Y7ubFS
cLZ0Z0gV3PlgfH4G1j7FwXjUUmSBXOFo/mLcQ4AUSAjzpKywP+IBwPzZxr0dSEwv4gVML8POD4NO
vL9+2wvc6la7vM8oOh1BqBuBT5n5jLogm0LhqK/FhlkcrI1iw5buEd6QWmF+YG42qLbdT3Fq21zH
fbk+a4lhQP8JuFzNso9kyZJKOcMZvHQF47hbD1I0gQ3tnrY7EYSiOZtAOsntamx20RNJ1ckU0Mt4
wC+2Bso006H+8aGBLXSc+FkagM3P0bpwNlHn2EcxcPN1ucgxjlGD4rxdfFhhytjpALvVs4GjkLdH
0hm+duI27SBIUC+FDSkchPXAoml5kxnzMJeGfEA8v2JKKgxNpq1MCZbP5vgY66IbOaWNagSUHO61
pRkN8kYa4E7iwqVDgmab4VeCUOGxVaWpcD0Z2Bj32duV+tfq2H2qGFRrGByD+a8vu06baETQLnvM
B7nr7sxvhq8iAk+DVstX25OkG6nuv6bH5eu4sNusg8+fzn+MK46xvNJ4oFKycjJb8tsth/MBKQkA
v0Yjtmbj7ePJoXdd72ScGRS5briCZ0XuWP9g3pWrErcxyp96/s9VxsFbl2xb/K9BQSy1iRtubvFb
yO7Z/lA6Xd/eIBsFNMRbMrjxnrCLLH67Ca44lqPyGojHYwIglvyCOJk3EHleMtneAR/BV9htt/za
kyjs/j5lf76D8pHSBpsao3U67i1UM8l+/OixMhxeTTpLN9p7RdIVopkYnDMNu/wASsluQKiY4NhG
Rc+D3c+5nftGFoW7IMg33OvzoGberW3zBqEr+THGK/Fe8KgLKJq2EvO1fOCJnrZ3o4pM7cqAYFue
xEwshd3rO6/D7KjMI3Saa3LG2FKypwlU0Nmf1RX592+eF+OlWaGm0GE3op9VY6ifUoGu3DJOB2Ue
3Hb/Q5drM0Qe151VM30GZkK9oN32NQYDf+e7irn3VO/uXVEKJKaa5A02c7kbvPpXJGhg6njtlhYf
fn1ppR5PY2p5cGs1HH7dG8HBnlraOCpvzTs5VfEw9FLsEfzGnhza5QCHl37ageBe43ONrHbh9sHX
deroCc/7HHH9RqGcLP0o3qtkpoA4pFQCNBpcWRQY6+7C4b4jtAyWiqSWYYmKU6CB9jN9OgxJUD5r
Cncx25WmEt29pri9JA0taf0H4AAUKypi8CE5bp2q1SfboH0gJkHWFp14tYQqmQ8lUVY3EZB1q+1T
+1uESaywLfGWKxi+5aLJ5u7UfRhVs3QPJH2DMUTxUC3IFfLMYsOEDZ2CCE0bqPk8g4f8/JCkYwa5
U3cOSeXFGPQwK/aQ7bp9A79bKGEM+dLfgMjqCCHbIBc2vvlEHtNvc0nhGnxIwh+Wwwd5qELAlhKV
V6sdPxhyAZ0xiJAUr/9HJl6w32GPmVWVtPLUfJ8o6rVfHT52QFmh5Rid5njs6ylLEghKC4FmzR8C
YkUjzPZTOMAwltf61w5fxJlMI+/7R8rBWL1624NuFDqX4GvT28kLu0MnVs/XNK6+xv55/BQ5a6iW
pbyYTaOoFdYjgDOkRplBi6G7SYXGVE0r3fRqHmbqAH/SsbfLLO75/wGD+e1zmfZdECMLNew6H5G2
0szGA6PeQF7h3Of+aHGn0ei2H6Oic0vZ5j7pCXgSY9BCbu1qjJ6uyoOXlJRmRL83BGTKPQeJzVLD
6zPxHP843fFXGhSVou3T/eCARtk/A0whS/NGpdUfIzOT+/da4adMxc0GiNm7KkTFk+QAm3u8yzXl
oqJm4xq5K9GQ4id4DJ9dUEqFVVwozhPGcIb6tI2okVlIeUI2PRWvwuRyP8C3qD3zM2K6+9W2qF2R
GPeVCcz0lEbjFd4QPT5DwLmIUHRJ8efgAt6sbVk8XtDhRfF2ltMID/ZQIFLv+jT9VVLngB1cHvc6
YhEGfIy3M/gTGP3pdXBOfB8aCyreGZzZ4xvMwgs88E2FyGXPRmk0nMYAnmQnNrpiIHoBP6VkrCK1
Z/btwo7HT7xXLqquu5nbzLTZOHfa4ORGeZ0EN9FzKTtEQwitErejLWJg0YhiJHYxhWKxL1XDGWZ2
tjJpvLUn3XSs7Ki4nwpKwjlq2v3L50i3V/bQIOdindC8WjQ11QeSk+NiJu71rmwzSGBJw8vHtHt6
D+U5PI9PWqrsR1AN6Fo4DI7xZ12oDwtPwXmYWM2POFittfMj+biqr/uTXm5NJcx8vCw3lngTo9wu
HX2BlAcH3PNmpyph05gd+8omSRSZHtFWZJpAj8dXNcH+KRiDUO1RzyElmfmqKICbYXCXHR9RapNq
CT9zQAKw/LBindSBvW9ok2BFEhPKUqgk/U7vJRxYkmGDfgZUTRgz6HQnQlCWBJrpKC1gBiwAOpaB
gXYJKaZxb45FljlKa8pS7a7Pb8wOzuPgUXgEl3s7rex3wOW8dbvL3b3OxshR1fUA7TJICxS0H/Pl
vmMYJfwu2p05miQ3QO5hT3rWsrk4AOSr/lCCmBbmbzKAZVxRor/u1DWWrbVihWTk+za+kw9hzSOH
6LU0EH4BVW6HEtfw8+m7SZHFOYTPvmlbd/EKQxqVXw1Q3JE8gIduzGQh2RNPR+h+h2l+zvI7NkiS
Zg8Xe2D/GSmYRkiYh8UaEEnjyLdmR46ICulArey2WGpit3Yyaa5JpAS4ap9kMWhccDHcWU5Ad7IQ
bb83ol/hU4QdAk7uf67meMlGYxbvAPDdi1QE6Q65HFm7ky4bzzBUXqA/JNkAujuonJqSGAQCnvHE
mpQilX3x3C+1b7GtBkbcW+01HBZWqnaHwiwMVbwEOl17oIj441WJRzpIlBF5DciwJkkFGONnQSpj
crEDXDS/6I9TzyvbrNS4tAwXTUInj2s0TEMTqnkjud492BFldhKlqlMCtQekl3XCMZxT9sjGHqaO
NMp4FrHanLkOolsegdDJUMal02ncmSILNnVqdGeAM/ejGMB6zxUDTYrkAnNuP9SAv7I25abS+0EU
UtlL4bkHcUzsQp3CGTslKyOQ+ITEgFET+zf/WK2/2icmyxgUbDWagbVqtScaDE7Nfv99PfAkH/Ht
lYrBxkKxZ+pVM1umnt3y7nQOiCGz8dSWGkIgddeMhEGaT5t3cSwQlax8VByrnOLLGOp20rgBgipz
NYROyvqeTYKBGONY+QYtzy4dVFDKkaINVzoBqFcDWAOGi7GOQLq2aEOowtbHtQhi9kPIh520wh6t
obid7E4gP1dc006XAaIKTeuSaN+ptKqfD+Z+Fv7khmUR6bTUyS3UmZvPySEAe5fm2mR1Vu/l7ti0
uJ7DAekQ7+snMXEjguix1fiEeA6Xsy/xWGmYMbayDlmMBVu/+0cb1S6QbjKVtgUQZWPWgApIdsXJ
hikf23xzxrxbgS54nstq7V1w74pWSAoefu5sVdeWL1vb/VvcdP+uN1JYz0Lt5OTy7QNn8rcouhP/
LeKReoHaIuPowvKAwyAlK3IyCdNbUObl7cCNKA0xmCoCwYMOjHThBWYduMpYhEQse7aVSA30OrKQ
epzMDK8On1YEUGuvpQPm2DtcBZs2bxF8Y8FdJnnyhTlF9xDbUny22JIllLiz4/sgcQjYzTWYFTQq
4E7hzBmRNgksfJQPekzpIBQKKCMFOCZnQkuxP5baQ2Gb3vqZBIXtnhckLaUEp5ycQ7OOPy4oEdiA
d1L/hpl7AFtTr+AcOH4k/+0ygL9k9hN1qFYLycthKecyaPfhLmgWi3XCz9o0dpoRIRvrQaLkS0ig
FrA3FIfcQls7MUtzxrkzEiSwYsXuZnuLpGkvYijdSeLD98JU2Pu7AQOO/2D737orpK3EXDCQDeoT
418NUb72b9qKHoWKal634zvtUJ4URvE5bWAw3DzwO75vxyiMfw7XDplWh6uSrlBt69d30eny7dBU
w7BnGveNyBUU+yfz/SAWsdFoGMnZR512OkeKWH5bWy6xC4kXpAJBrLOmxHA+0szq0Tjyn+IBGLSf
x2ZVqHVDK2NDA7u/CxWTVHXzlXB+L6mbcM+KvzF4s9BUjntJ7EhiU2glqR/BSUaiav2+oaU/5seb
0SD3ZGwAHiK4hQ7qF92HBNcCL/v+WW7YeorQfh5IF8ZU+EG2OvyF9GsyqNdO+3/KGmOb3Ps7qVs8
RWsRbhY4ywWYdoqLVYwf5FehcaovANd1CcDKVGYOj1dIZ76lLngRgMKB2TzV+EgQ7XTehgUoKcXl
bVn+LxlERvmeZgLSTDQNWvxTiw+9yrXEPeVon1O4mKSm2kVEvc1/qbGGrWLR92MsIcC83Bbc3kTr
YJhuCZRTTZqsJj0yEHYKqWuXUH9IbfSbCgiL5/uKSlLQhRnuJF1RfIn+oe2clyaekhCSoPpEueUI
QGbhn+/e78s8tXUSbxpoktjF0NWso5hxe7wExS/O/8NkewFocCTN98I7bfH4spIbXBKWx0TzZIbq
YroX2Kmr1rxHeBIo2vZPHxvYEQyE6IGNHviSkQs+l5m/kpC9WqGMs6BCH8WHa14VEuZjM6k6p+tG
zSjwUzrQpDbYu/u8OsGUjaJM+N4M4X8yBmkpprOoQwsym92WjLxQ6jmlY/qXNzg1T3JbTYWk7xeG
+JJRzuYuL87RIPEciQALgpSb6HSguUD2TYPbLpBS66Yb7rgB1A/unUCc/ygjsppN27wKwr9K/Mk2
vWsoAcCLIVmPyXhHfUK/qXQ1dLPRLscEycI4az9F38e6dWICkpR+52ecksb5ZbViZo9RvXq70HyY
U9G4+Yo2mJdIvZrD8oS1eS5KxAVdeRahCfegC57mASkQ8pBg6Fl8ZfalPVTtQl8PlfaV+T6snDcA
+dCDOThBUmdQ5Svb71RnbZe7Pcn64brZJCoCIEtnZJDujxgtLSYiAzSN5foxztwCOqWQmsypIgJ8
zfvxPNC6f91hePabnZ+FEQaNu5QRVbd3m5VfsrpOEWJ5566hPQ5DIGsfnvGgmYVZcZmrr8e/yN/V
IyuvkGRa6zW0CU6MTY8JW/lLGrEkpjaegmZwlkezc9GVpWBmHuzGIMlNP//04/keRc4Jiq+3r/M9
jDj2mZaHST3E3d5lsri2LG2NNiOcUZ0qwM1VdH0e2jdEtgApe/mBlZkWpKa62brWF50pexq2L0eY
sOW3dDm5/z8EUIQoOcnzOzOtfbrMZE7XEjO5xiYoSL6oh05NDCPHrxTrjJsuZX3PhSHsijWtPIep
bUtLBY3why1msw5+RlVa5zQljiAcnDowv8H5x1o86rhx2bgRO17Eq9UJ2kS/WW1nLDNqG7VZmO5H
N55B8FEvB9/+igh+mU9GzKg+7wdX6bLbR0zU8UNwVWRbdaBVBZNhHlDhpY2yT/qpajy/ZZdkYfHW
u9VpTWKBzWhr1FJdra2fkfBwlleYS4z9blgyMrfAVF7fFSrbsQXJX3U+NlizptuHHoib6VIpwP9J
TBLLgzuZgGEnYd8y8T9MZcz9fRVAPuX6izSXyB45OcB0iwFQ1E1tAZqttVJWI1r1Y3TI7xqsM2nM
fsuXBgGZI6deM7OD0QuQq3wcqaho3ndYcvra4+tAugmmJ5JPgaG5H9AyYUIRC9PJ+wouI/aEMrdt
977OKXD3v6Ptqy2r5+Be+dmw9Xsm+P88rY44RtM7eeK6u05cLk1Dvpw3m4cmAngQK22ynskEoiAq
6wQ7hDCGF0VCXFoeEi82uXOsb4ZfyVPiZi9/wLDksxtLMnpYaq6csSq6EeDO+gebemrt+lhkul5Z
k9frFQl7hq41REJKmH/zd8mh36DyS8KoHojPJr4/5YCgb1w7Pf1WVOxZu8DqX+TD+WnzfJ3EvB68
kcBc1u5SIUymocOwUxL0F9Ef70E6BuFf/Oskm1y+jsFCOY0s89LPlQa6Bls9i7BrGWwqV6VKsCAW
D/hwHlVKnldcWFtxoM/h0HHe+LNlfCWj3SxcrO7VGDY1UFCGc8S5+GQY8JCxa4Z4xN/5WFeEFslM
Ei5C1ukerL3njtsV3i1alPrXphmvsrpf6Au3d7Dh0jQuIL1T5Ak3EvyJoJktLljU9a6durIwsmff
b8jQVwdqHiyS/QXcSe3aNfc3UcpJg6Bt4DOAYQD2Tqqmyso5FA2XIXcbP57wG+aiuQr9Q5Ia+tjr
ykwbgeu0cNCmeV5fZswR5rjgVaKf1WlSU+jSiOzLTb8sjK5WihAprCjps3KDpYcY3g5rQ10JJnqV
1DtKNtkRENv68GsN8dj+EEWnkTXeqa1RwDBvttdhhNRwDTL4meNlK3yZSkj0X/qe5vBX6mNUNblc
Uvv37QnK91oW8oVDP86o1msMGJ+jJe8GpSwjIqZDbf4lO57K8PcZYgfpVW0gO8TwSEX3LCu91tZL
1pxPyxxBw1iId9vrKuz+e4BQLd8KP2Lkl1jVlt51hQOsRrt+vIFOwFFr2J4zLJrB/+pgrnca77Zo
OmB355gsnSh2UyRgnWPWHtkLzSjjGKvoi9oD0ZkSjtsZ5SuHpNa8rmVsM2N1SOsB0Br6yy2IQRfx
g3Kfq23H5jb5IeR3e/ljKCXdzza3oNZ1/jrYR8GCsVyke4ehswVSO8QkeehhCV1GTfIX5yPCRQUV
O2uc/OSW8EhUbjvVU/0IeosljXBgBgNVFoVaAFdFYJgyjlyKMYNMw+uaVTJJXfWHO4qClMWDP2dZ
KFXJfkLE+XxJBWV27mrVgXK8y8Xf12Fl9FkktCmZrWoFD6ETqf/n7kfn6MnU9aV1R7J5mUGC9LRV
sbeDXAfvACswn27ODnETIHwNxTnsvmeF2UA/d34R3wkNSd5eA0JRi2HMby9RnSWDDFw5VshnyYQR
NfRpsYNkGfe4WNR2268a8RkEbsYPvU1FXI6eN2haiB+JRk0vv8a2uCvT878yzypAyu7JNpWPW0Kb
PsnlXmgQAkdGDfRo7cGa91hWTOzZgCzgTHyU5v8/OXcSV+7+HBYDYTWPAvFPwpdl7mvXNIoYZsha
jZfVZpsr7HnZnF7bRAWSny/2waC+NxsbeosGck5x5GuKwCQOWncXPZDeY9UeAsOV8yNrZrIsRvFX
77zQDhYXCTUbq+fGonp1s0r30reDF8FC4T6rydztiuzLL5Mka3Lgg5stqCaxVUaM2m+1PO9VaIUl
ZSjtZgxKOZZFI1rRVBfWGLcePpRhwEHuG9gZ9yD26WLoVlf1IZiWHZ/ZCY4ayMDQqPb83NFxL0Xh
0Zet2P5l9YIXRa+Fnh+bV/6+LxtfQV2noRvo7ieLw9QMgArJJzIpxWaloIJdpKapTVMFTJwxo9uQ
RvE3VIvLoPLbD7Czhx9C0us9ISjdD6zGSC8ppxZL9OksiqShdCJ0XfTNRhk7iklHJ8KHivi0hwwd
i+vQCjn9tpgcWQfgKFHJZYEqR7w4UIY2QW/FCiW2Yy1ecGjlBoEZKSrg0jVcOJf8KgHhq7ubIg+X
4msicPvVB6W7VhYvRzIrgmdTrOsWKe0yg9QcnthGghkJ3yDivizPDxIdyVBoOr15G1+CwyPXmXVW
DkL3ZvS4f8GNdYNCetCiiY4B2BVaheLxbz5SNuSib8AjWlwchdb4OLBXIsUhlAs10s1/8qjlOkgN
KsvAFXAnNAioQrJSETs/1l4U51MmI+LC9pKAHSn4lGORnDvCEqMDdiGdxebqnUl6fEjQcI0cILaH
Em2W5zlvgDIoan9SDwd1XgjCgARPe3sgvHyi91b0T9NultctexDbBJLWK5Bj7WVTR2OOH9L/cTzX
3ldJBVBDr0POX/u4glFrQKpxydOo73tJ5N5xeTPxgi0T8UfQU6RaVorWbLK6O3aoYYnwJjPH/F69
+uEZipDrDA8xYM7ptematERIe834xD9H8Ukqdo7kU4cnLqndVpqOyjTDo8a+bwuvWLR6Qzrq5b3Y
hr7jBG/2+/AeaFLkVLCCzov/jQMFXGrbdQhhYpSR+3Rn3y+O3kBMO6zvNh3TmlYarqhi+FAi/vxq
o52PcaRdmfiUp0Ohpr09tqNJXXrWIQT/0Q32m0G1MtX9DCiSQzqPJ9kauO+AUILDJ9i4muzrLMIP
SAdmpBnOupExnOZm/Z4VRJaKUEK62BAiuOdlEtYOAQZffDDmZElPmhzmIlo7xIQIPUGjuMQHKZbR
NRLyB9OsO9Jm/AIS0EnxPSOD3uLfl2HT44hSQbsdButFRiFPuZxlxlBhPzaI15s/IypnYBDhur3D
DDsXugpEl70xFSm3icIbXpxoteVpqxZF26do6JuUiQ1zCU91KbHWX41dQe6xQ0BuyRjS7i4PP4WA
hQfhwEWTVlDVqqVfJU9xYrTdSndj7wtfcU61LTf6zrGqBNfoKUMOqqVRNj3Sm2UuOjFhAEAuj1cj
1GINLw1yh3OQm9hsG4tw964V3Xytgf14G0pnbnokX/VWkvJSt3Koq8+r0YV3uGPOOVweK5zo0Wop
pJhtPIEmdW385Z0OMg3gC7Xm94BMepp8rlu06UFfOdrGESfiqxDTPlNPbglhydRS17zBvbul4D5X
YOdpovk9bbennon2SkepaqXEzOBnx9muoUsHp8X1lzXTuGnxzvXbYfm5YgUwrUSHmBZIwZ/+vGTu
pyw9WBg2ysTJIdTbeEYWDODTX11dQgDSZMdHGhbPJ5WZUFv5AYPutTep5MQK6lj3MSt5LQVBCJTB
7PMFo58FKdVGyB/n1tUCp3gUVwe02bHd8wRI0HH3l8F+ZKnjuhspY2TfUUmWvqkRux/0yHPJu0X6
knnGE/feDxU7z3LHQEzft6z2pS1aJP4iqub6hNv6vvyRSDPWr0v8+OlELbW78Rwt6YSYc0cG/Ahm
/kB71PE09dMRrc90SI5eRImbBRMBHAWbh6j3f6JeZPlhBsiZYPZtyrWk3M3AkG6wTQOBa/ttsnSn
PKqIWJzo4iVa94ulddkJg8K0B418bxw3KGfG6UqKpxToza4g3+uCZa/EhzHZAyIu2DIC9eusgOaj
g1F0PcAMExuwVUstV9Y9+I4FlbQRgoSCgILQw1zhrTr8gv2y2CKA3Vq7Hx5J0yHO3rLM3WPT+z4g
oqNoXs75tdD6UFwiY96MslzFP7od56ZJspeogBT9K8+WPOhj003DRiRgC5cKf3gnkD36mGHAOHdp
QbfP6IJbQuFRCs6GBRKTxWUsS3+RYppvtuKDTAHfV9VBqk20+tLqmokAV3r/bGpvT5X4HmVkxooB
x2qGmTPKR4uuV0ITtApn2jn5qZ3P7B48Y2YUuhvD0QWukC2trWNtwNnYuw8XBGcSLfubKW6zeueH
PCO/V8car4VNfpZq1u/1vXdF7rYe9Li5WJP4rz8xZzoKgE41GqMb3hgKbM1Dy8NoLYrCHASxE6Ao
+FAjpadQ7CXnPgyco1c/HPztGzPZY7MJGN/IN5daoqV32Sx2N2vs+iw0+dMK3wbH9ikGk2Ql4G/b
AMA8q5KJmpkyj6321T/L0tRlbd/0ZCtSxJ2Z0e4MFo3GxCUGw/Q/qB9mEoDzTEj6REwmE4w9+UmK
L9wL2pGIDz4xUnCv0oEw+9F4gl4cebuJl79tXFlM4/9esfaNIWn0kYVNmKmU02ZBuya1V7inCZXl
jeZCLgCHyuY2dkbcpX9wszKg6RW+opm1wRsetQOI7Zwu4+CpuwsCjCJglvRQCSLEbGiTnZeFqvd+
T8AYje4VbIAMNgEDtj8IYpsXAzlme54hAQivrRSYVwaX3tKhYO1ZAX7kmv90a0c82RTw4CUPu0fh
pYbeyVB41fPk+SARcsczGYI+XocZ/w4ER8R8anr03bIqPI9cxNmgOybiOg6tYzledNJVpKQkz8m6
GofsyRnK1d7gg45dqakqVsAB5XIe/vvk+uJyGXO8cK3v8s1j76IxJyHiqDkCepHPvjP7OemPJjT5
+8vMGgDwRUuNsHh4mw9uSTEEiWUzn1HIfdDD2J3jx1sMZvf1I71YXw+/d+76Kr86ZcJ5R0nTAsFA
nl8WCe+xc5frF3XGWoX9zFmEQnFEmhXjkGljEvMSmwtpq0lY+jxSUSANJjcfRSqdO1FxxIgouQZR
z9EI53PwEVhXfOzEX24CeRAbHi5Zi7KKkUVt59MFG/RmV+RNem04ge5HCLQk7XHM4UMdL4Ei8az7
uoeSiw1aFOICvIF4SoPeGY9+d+hwLs22onslz1llD6QH6GJ5w0f82ye+yBn7QiSTE4wM/hOauQP/
P1nwqXfy3PCmAVl5i/9t1+X2ZYBI8ztPHaMiMy0CNmYXod+hS6gUcC2fmbpCVaOCLRp9S350XkGO
Eqer73JzeAurylbg3LL0zXlTCTNGX7sOhVWOBqHGjKV8CV8mWAGoQVJKDqWgOyLECzOO86BLPt45
+T/K8PKkA8GfYqicxhMSQ8G8eZIkTIBxHVtfrtlcoe/go4368jgiWB/OXLvSq2eRQpCp7qbVnEln
IxyS28Riq6fXGkmV+Az93A3mcc+rfe/rYXgjJ2GVRRHPJQMGqbBfMWL6OK/K0hHU9BMRWn3VoJn6
Tgjy2mEVt2TSPEHp4oyLGls7YlkuigN1mLuDVc8PhjYqv0e3k7+jLi6ytulR/M8oByHG17Z4ecSL
FxtsmpgY3CQg1EzAkbz6BhjZLHQnWltnXuxxgJpVEpYCajaYb85AL0X79xYUvwPRb+9RFhATQKYQ
LZ+5Rgt+H/YtsSSi1YL18qhOX7LI4i5Is0Ts1s0Ebv9ezBSuT5JSe7xfAjMB7XOGXMcOtgdMZEdZ
7sudUDauC9y7IBcgA8ahVUWh225nYoTveZEtGIlLvqqjk5OjIoeCSnaWLy9KsryJdBIFDxiI2+2c
TUGpV5vAj9qCKjbpLElyhIlShCZYs1huGa8eIl/b4tftqa0ldwmXlUW+0CtN25H8ps5PsL59ffIq
uac1927TUY3UVZ0/GzVJIYbu+DEko+u4SghCDfP9r43/QHl9VNeliVuawRRlX3h5cOaJeaSZUmea
oa3pMsW8GW3TmT+vkRBRT7aAJwWqwMsyisQt76/WuCreLclQLF5OYVBAQqN68LyNeDWOi1Inuz7v
d1iIIFekTrEDTr1nqGeeZmDix2YCTqswfOkq54qVGWXsqwuNZMW2xaN3V0Y7KQhR37Ia1KEsIEVN
IGSuNwFXNaDRYnCKqySRalJD/QHKgmEEQtX9ZMDQChrUeSLQl8qpjqCd/1KIwFB3P2lCp/kW3qOo
QrYD3RysMu6+bHG3vso4XICdGzHkAVlM4mGHT2abAObD0KlIqLIkK3sSrHTqfDegnHBuOkKjYqnV
6dC/o8BnCmV8AY219kIqa+fs4Au1b2qZS90VqJac3ZsrRmVCNek4LGuIWWrMZoZwe3OEAt2ySgsV
99jdqFePZHPgZ+5ZRmwV8BM/jAflWa9PlbRZSP93u5ZTwEguK8v8oYLZpkAWk6h6yIYmho7KHSh6
F926ESz7GIXk4xjNJ/GURQ1RhCI55xr5izPcaQ3xnQJVkNAFszmrp+aYKodf2vWW4UM5ABXscNOq
V1nDntfp2F9okFMXy8jcSez5Wc8HVTnA9PpnR9FgDYCylfIPoCfSVPhv01EjevDTCGiRqoIPhmK5
bAXrT/47YdXyyThclF/c+VQmDfOlSOzuU9YAo8ANhtxhEhIQorA6oQfVJvY6wxUsCC//kO6PK/XP
a3uqNnX34HqpHaLFTTLxDL4ArX8/qmBwLXQmxEegJ73aFTRrB6AoR9r2iJ2RA6vayhX/nOXlbWIh
ozFxcMZ0nrvKnYgw61Z2V3H0mqkfCilQTSXKohbOh9NBZcUv6TwhMn7r18fxeGSjGw4CyER/tYxO
2QGRe8Mru9inm5NA+r4tRoxRUy5PxazrDbpWmoPnSmzGojMm4b0535ZaZmnDnPYc66Y0T0PN8370
P+Yiht/K68LifFfY6XGbXvg1GggfKP8DqOLbj+Q2NcWPlVt8b8TjjEMSLC621n4Ha/6J7LZKs28F
uU5BLouZTb3+wZeXgIE/FTE1wgyx0Z+BYWQrnCgMdJEJu8loTKS5vdAKQjw+7d+vpviXEvrCnplK
4zj26olsW4eMlr4rvUAE7HanNK/29bIWrlzDNpaRH1GzfZzb1rmuL2bvk9u5NC9/710gTjRLgS4B
Luj+JHlb9hn9T6XgfC/FzdyjYzplBmARU6epsHeCoLz7bduOCyOdxs9TVhQb8IUfTyJNW0px9v0t
21e2mue3CnyKn3GB3C9VJ0zUWA135AjLn5mPEQyr0U+sQqpZDXbv78o827w33Ub9oPYK0H8QUyxz
jldcSOotWMjPlVAT6SDU23q9XkpLG0iCQ3rKGSS61TsZs9sL0NZsaHdi64unzJhGtGwwc6VfrMxG
rMBbH8PdLgdnXaDLzaArEezzL3j9Z9GHBz33qFxU7pKSFX0lx6BRg9mjZp2KMAGlyXAOC6p092QY
e1m4k1J2Fu0S+lYH1YGyuhEbWZFg1EvFnETA3cVcnQVRutdbVbQVWioWx/h5AQBYzL3UBXDxv3IW
l+WwsHc3q01XZqnsYB6Gunic5D039UNyYFwLcV2rmaqYO8+vUNSP+nW9zirt3ZSITToE7nqSd3Me
+kFJcMQ2spjf00RgrhfxDAJ6keRiNBQrLDMe1mD6/1Rxv5w91l/dYVPgS9tnqMTpFjXaN06lzIVW
KYXwluLbldyJrreJY6IcPsw/MiZX3Vt5WygjNktXjjf78IULsIwBkhVtasiMexdUDcC69S+DLWmm
VTy4L7JX0tXcPS9usBjr445X7fijA8HQUaKco3UrIvtYvxoWFaC7/tCUvfNqgLR1wJKnU/S4BoJ4
+TKRsr2naowcvkEGAnD9OSxOkD9iVmqFEgbzh7NDwGkOYCzGLUoJQ0z/WLNwHEpCGcsxn/aLrKva
XVyoJsHDGr8kYYnZi6gdPy/kOxlo0QIh7qhmt5EUtgJdS3QAbqXqguhi2K2dScj4eBGdogRobRmX
yluZtWitZkLlxrfpM8F8u0rzGhT4S/H1eGaZ5ThiVC2tEuN+N9yLUT0mpjfUEyu+LmVUImkGhDGa
T8wFzWbzG1tw10nABs3MJLCRkoRPc21+qQXr6F1rs/BlHeTNNDgc0Uz1pEN3ENF6xKPOmzxpOgq9
twhmiJsXPnCfTO78mCnmXQIrykRsCDlC7v1pIOhW/1/FdqsHtVTswMcv4aPWWhn4wx7CWjYDgObw
U8rlV3rR2y8csAhdrspTWrpttOdbfHS70KLDQ2jrJ9KvAWEDjYE/8AZM95Liov2sx9L+PsQxODqC
55SkfgXoz3F3mo1q8DPImwUNirIO8C8YmGfPBfDmjfyvYq3UdNnR+h5bznsNGi0srnYicWRDJ3hK
mUvFbBw3inLrUZYEhuTuOv1nEI3amJhDLjiwxCtE536USywYcTGQnvU3s2GqgOXx9xPdXDuc9P7Q
HzMiDXFP3Cm/vrkH1R5CBrdUVx729KipE5vZzrWRUpAyNhdQmmBATvK3LQBm9N96vzjf3EZfqQv2
fkqwfYzPOsoaGwsGNZ/dw1TByFEE+h5g0SeWiRT3h0IFXskwM0ypxFKAILckAjZ1EkUSc7dlJx0v
O+JFP9603hjMnx2kp4LHVhakZLwzG6UaXYcMZP+KvWU/BsdgDK48Z+sH4xq0/V7hpLQ2md3tlsG4
1C+QN1SCmYI8OkrIrIc62bWGaXNleJEcK1QZKpkYhpEP1X8GF4uv6SJoEeB45BiyPWYxjUz51vFj
E4Sul7suXZQXpBwl2jUcmyOTky86CwaU/HVoUYR7MQDWFdNK78RBZYcWxxSqNdWnXspj02+eR89K
p8zycLLm+7VpjTlc5kladOk/cnjL8d/Z9eZ72P6ir64Dx6hxuB8pmiXZwjpaW8RjqA48gyrudb1F
eKJJFtslGHiWv9Or4XAHmR+vQKL6nuL057wzZu2n0gZ7KTkEmRbjGFphc/kXizu64o6Xhexc05OI
Blh3uVoY80mSGXHQB9JbTAMJLrU30fZH7ujDoHwzftgekHqZfCA4ErY8zFgk4iQlZDh0PHMrC67F
q19yuc61xZOowMfjF7sH7AxbkOn1k91PgzFGxsY5ioaMNM1WLIgvy+fZCoz371J4H4J6MLoEZx3j
4tb02FrpC0Ypt0bUtFMlEhjk42cjqAuioqPcUxqTvAC/LJDAO2mJ4aUPSOXsZudc3vVe7VY1pmAH
VKAqFNys1dhdUmd+TtmuiBHPKfOLu9rb9V2XSx/dpqGw+PU3aq604i5U2FQIi6Xn8cqb2zz62X2U
E0uqaanWI8V5WL+MGPC+IghfftVjLfNRTyT6uZ4f/VgFGndOPWISrPtrpAXMgu5J4QtBdplPs+u8
khDb3U14CpCV/eHx7Qe2jEMWFrB1cyvSsDCll769Zo6OQTLidJsyy3iSNLgOjA2FjTiJO9QAUgWa
k5adUH2pAvkj+vAn0A6SnnfmeOt96s6B+kbfNx11+5zZdzKaYtClMyGHJtacX54zQvisxY1eYYaX
c9qgBwIBF5K4QS5Wouw7Knyjwdt426jjKHiAwWn1RuLMJYW/TpG9k4JPMz2jEctw50BAHeUZajVX
pPNBhsAHGyA8cqCti4L5Zp+ZH5wyhmnsNgwTSxZdyXPnzJoE1Mz5IftQ9nTfOUwNBXu6Cf6Ij71P
4RPmtH9jyJt7xEqJBxXjjpovtYRD+c99wuWgjxaYc8KSLhjJt+QS30Fbm0PtC7y25lWnujq3dYVi
XpYAETRP/1Nc5vvbJ7nLsOYd7G9c1dbud8LPDeoMPkuZwD6zE3XWhGjTKgDW/bwiZ4vOMAGFyLxd
mP8IRrxiOfNWeV4C0OC6pnwhSM/Reu/wBu9khu4E8bGEgzzBR+g7pjHygMpJFU2mzc1xadfxKsh0
VmZmSTmlKHiIllyAdg9lV35MeZ1gHyOQO///+9wj+9oEET7wc8Euxod96a0siAKJsZyQeIQxxR14
2UYVHzH/VBvCCMDWhstm+I2n0v5YvRKYg7koVU0E95xOyH5MsSJQXLvXksxLAkKdiT7gNW6oLKvi
tgBnzKDKmco+ozLG4VenTPpr9OX2iIv2Hq5masp/Qjlqiv9ICHxf2rxDFp6lVeCJWBkLqpWn9gv0
YZNdCIiUaFzz2gWkjvVCDGpispC7jHqxfLBQTqahFptWW+m1mx3ULynzBFKu94XRN9Nl3WXfYkKN
e0cvJP048yYv+H2ZjHWQg44LDwv+WnRFxgfU5LNtGfySYmzQVBx7H/Stwi8YtqCcBqLkBPyAEc0K
GVZiscpmy4+KWo43lyM9yHRxeBxkl5g/zpW3NKn6svJodasyzeyBgGWtxoPLXgPp+q9B/zq2lX9u
FcjMZb+qj2BGhgUVMxZd6kdLM+7yHUTdlUYlj+djtmRUhb8qKAehA230yFdADyDd6B6hD6DLN0nS
zTow48927vpHNsdppmnrsN2HBMD22Nc2DgPwANuJGrc/wxlwbEWqrkSMZnRs6bi1XyKfdvijjSOx
DojYFXU603n0k90GkTSYTsQnlC2e5S9S70CIp/f5gCBRwCKl2YRhyPpmDrZy13qU7ES80h0LRM0n
RG0GZ3O4xJZSIzFGe+ssg1lXaXccXuygru1MxHf6aatSDqXQiKNTu8hkyImAOrPPEhDzd9sZc6Ie
e+scLWEbinhiD5QANTJkBMmxjz9n+vJvQ3KKYz0AErTpJy5ky3gBSH7cRjlFo+4g1/9+KgJb6C+/
xijAhbL0PVbnbaIQCWKl9iwps+q4y/ocFwDMETQQ71EHP42GDN0xIOPgVU7GY2pcVdKCw4lOeU25
QHRY8FkLUj83M+fy8tKBWe3rQLh0lOhYbkAdGFwldlDUSYP4I+PgRWstsEAywQ8E9z/uLwORi4vv
NbhzO/LBLkxBB+RwGg65vIcHyUh6oV/HBgVSCoypXChkLYWX89z57oBCI5X+dO5c2OUReBDv0OZq
p0QPKtiNSNN164yN26LV4rJYtq+CmBtSzG2PMdGMiXqjaE6Zfvrm9zbOKqRB2fS+5IEfKTxRXw9O
Hv68oAOTr4itIKDAZho65giR79lus9USbyEfTNuBBG32KEAVyVqn5JGB72iVX4CYBVrwL+7ipRjx
N7rDB9UmqJQZCyA40eofqOKxB/T6Kj7fwedQsFIO7X50JdfOt8DT8d036yjyJf5MBMd75bCxDzic
Cn1HajewBNZ9/i6gsYhhI4z5txxN/yWlm5R5n/KlFqVrFOKjRsG6Ot/2lgaamVocx+nLiZWKKz+L
BdxAwlxz1MBWuERW42R34c9eo/DO+pux2L58Im9e1KKXAir8dK87oeZ6WsBwJJ77DVEdbvWwiTa4
x/lUkrd7Xz/QlZhLv7nsTtjLJsJwxJPkNRV8UyZC4U6/BpTfezrWKwv12mX4MLsD1hE8GfTozeiB
9P/fpInQXxHZyNayb72s2vOoE2pIb5F05+FsQrarkEhCc9i3c2ubh/tG+oGAjBh1DVuA1AHTsVFH
YYReJq4QRDrpKdVpMrGd6Eq2IAhwbZij9toeHKuUYPvtZ1q0KUlhZio3LJZj0Wb6/zuphbJWyhkT
ev065efjSRs3PB5fKZfWgSRuSf3x5eDHj0ZI/LRJEfM2eKa9vkLpf1HdJ8nTSjiRqc7COFMQmpsD
RmB4CYGX2kFO3IB9B9GW3OKeFpxtKM/HQ7TXLIIBhKzj5JOB4aAc3uLjbmkYt8C0pjp1s8Qn94VM
nOIGEWc/TfWzt/ilGC0JmiI4yB2//XaGaWin8vlKN6miKarTm4zDcRfx3ig0ChKyYVQgojtERe4d
drKipsxeweAgSB6g394pmToaCJWC0BRsv1O1WI7At0hn9bhLHsHY5R2poUN295FYPxtjmMw7eZaA
SPeopSAR1bEePChoLwAQjznYyprp0003QqkHeeKL7/O9FExcW7Dq8tZdFoyhjYT7Xc5NDmAFaBXT
km7ADaZPB34XcWPS+fxQgoPb2KuHsXWol1/0FEI3MY3SsHxS7asqLxZak2+z8ifxlJ1TNBo4b5nh
j0zqCKcRMt1a7pjFOwGlsKUH1zIv42IvYU26i/jEY5ncZTRRB3LJkFENrIMxMbLl88dXcJarNxCF
+4AKwmX8jZjjarQ8u5GmLPEIq9KooHj0QuCXQaG5cgLhTB7oyhRAYU2/C61k6vqc3oZBbVRO9N0D
wDZNceuw9fDzTLVABnrHTNLxMLktJ7mqdTIoWYJiIoO3XxLAb23v8Ear2EN4LRSUBfWBylJXZM5h
mg6f9H86LCwrIl35MpU2lQOaBDJtG/HgHJ2tQu6D3QGhVJjkOINjErFH7yWg0Rf/70NrWV13HBbc
miOoxbhhGX3vxpsOeLhARlK4csP9g7fM8YSb5zcQhJuODPVRdwaI2bRyPyEyYGNKw4eRAX1Ud8V+
/daUFiYrCpOGAWQQzkshgFebven7mrbLvgEsoraxQk0/OzgaLfWoGc+2J1dv1kmMbVHT1+xWaUSN
LknvBOazLsNDXvMvzn7H7xs+ja2qBPIdkfZMEKtGS+/IVY3ZPI8bASLwEgyP3v3QQ7sLMVcrAgi6
5emIB1KeiN/CpvXL70IxbaIuV555eCLih277w2c73Bbq6yoqk2iLjNdxWZBC8ASF0GixgPa1Vn+a
Yp0cyKPccjf7DM9QWb3p6U9rP6VZ0qXio9sw7+lWzDtOl9UFcG6O3r3aT9ZTgxWqQlhYucvx5khf
YLKbHj+kHxabDT837qASAOX2tBxItHZ3VrGa2vPpR+91inqrUa9E1xHHlRUioDS7Z/3qCPowvsMH
E72/fjo/g+Zgx0OZ98b6Vy1tDG0PkgF9JPgDP814YQ9rqowCXzhn5fQ6XoIVvlHyWkhxnFkRARQE
ZLuxCNgbxV4oBJ+y008Fp+fs0qrC6lyM/jVzV3pZFX3zqTaH3kNtUcfC9d3dZUzk30dfKMO6fDKJ
5Ed7G8mNnUAlLm9U6YJRJGGdAcDKLj9UIb3hxDw0etonupIcHfcKPQz8mA492mY8aI0HivD5T9W7
0Fp2apGCj4BeFsQy4WB2p7RD1nnW3ssuiWNn7XE4bG5h+dpTBOaUsFBSRmKlMElCwlP5ALv8u/ak
vHXzGkslniMuf+GJQ4HZ6UoSETMV5792+l0XONGfw8I4u8nWW91OfEJkfmFXW/OXDUALhsv449no
U43s1+ia58JQbg85Bq4tdfzXt9j/K5FDrKHVfe57cq4xLjHQSVThl1V89box8FqipmW6o+Ef0pjw
jV1m7yezE7niCTpltJpJ4ShWQ1cE6wRAvMce98CHTDuZDfdptGiJ2GX1T3mD9l6VNBLDIrCsDhq0
oBsFTOoOnC65OCMgqRLU+PD2DzaC6iw0trpDWGGgN/M5zG0LglRAURs9tyXBwH3HawHru5S9NK05
+lzWUaUikJIL+7F3TU4bziQUPoCTr1AZcw5X/NBl0pgGIBHMnVlu7cCMwDvV4cQ7cPAQ858MgMDq
9hYEbKkmVc8+i2fo9pvW7SyafAw1O944wMeL3QEW6YdAJW9kwKwUpi28myDCqEiUoTr0WCbB1K00
fCDS5U9WeJBDMchuNNxym+gkxezeEuswqnEetX7mKTy4KDA6XtX52D1Le5kr9QQTzhwMcnpKRpjP
4Q3gYpW0OYH04oPwYJFPPyFVFKpXy5pk71zHS/pdjwEtsbiALcK8O0yHncFCGbaD3m78UuMVunIS
mF1ktAE03Bi0JOuuAitvsQXIQ/d/nGD/lcjtz64PCVAhqAEJ4dJx2ijEfdzOvuhMRtcqGf9G87Vl
rp7F/n1Z/DwNR2hxOsunY/izns6i2oe5HHJ4gSNRiqSURpegGZZsHljDFtQuO/Q3ANdRGN5jDA9M
RVDOU8LpsCPxDSFkyPV5gXETXNnNGbgznXcQ5kziCjhVB1teDg+3LHoqHSyFYrzh4AvsGqUGwWvX
xatLiUXCvGryEnozM5kSkAw592QeP+ya7zhypaI7/YSbDUk5nYT/EflL9yiCIcLvkCfvz5B0/cNN
cwFD3b30Pnf31WPCnUv2EqBzURmmpZcvv7dMuSWs41YDzA6bu+Tk6ZHzWX8Z/MlKV5nZDH/t75Vu
6LZ3Pl+LFl3WljuQHcardg02h9Lf7/1S8a8VPkH/hMHNuMq7fdCHjZpcx9y3tySya3IcU3OGuyyS
E7V/7Z5wfz8OKXaaaU7W07NFj+3Zcv90qopL3elk09gbJBITOv57PdFGI5X/yJ6W3qf8/dgFtqxT
b3bvonClVPfA1PIkUerH5xmc4mvYfozmdahufB7zxTC2dItKMcdegT1U+esXCAd+sDkXaHueOJQd
mhV2Rhtt9rwOgFyLs8RxxuqhIhVMCXSpwrhVJD36Dp24+db8KffaCrpJ1lJRnPmWLGaBQKWIpbaM
8QOEpL0D4UW+gpJf9TAwhzaVkJJyytCSwGSiJVByGSS9cSKsFTWkxgWv+/GZqFGZOFuzewjqsDt8
b83TFbfbB0aT71AmSYUkS/1xVP2SGpuYVz3tBBCyRmRzkQRrdyI3gdDBiXZduyf6dWAzEIcAY0j0
3s+8Ml6xRU/1n6xvT6Aem2TGxy/xXdkbm65NxdJnYmO8AMdk+Ud5Zx7/lers+VHdBV5wwmm0obmc
wnJLgEJEJTr63XSxFtrgUGGCAVs/amq+7DzWGib+dvDeYiKWIMkqFjUweKJxYXm9f5pD+FU//lM3
na8gC6fhWLO3d2GVq0/M6JlJhZRyPlttb1tPMG7fZ8UfaBBI8NlWZkUycquH9UJSvxILEDeXJdX5
fSgP/x/5oZc/4PtbJgH4bBur7gW0DwnbSdBPIvxXwTU52/3oj3Up0xXQ7PeqJ/hhN3qpVh0vVb5U
JLxSRnO68EbDsYdH+0Jh1qlirGzp7ea/rsAFxZYXLxak29AWRkxjpjVm1de3PuK/Gb7xiuofkB8M
N35M2/kLmEMHnapXv+U9YdJltVlUDOJc7F7chQ7UCo1FiajABE9COvcmSoQQ8AQVQ5L+AM6d3AA2
c1fuszV0QgbMpKV2ECyTxPB81tNCYJEBy6Que7FE+77mdJfRmcBdahaJjeH1KOEYUhcY00oBZUEc
WMTiaDO0cXaH8Ge+Pum7ue+ycMHObJEtXqhh5k4MWtAEBcWhK3xY33+0JgSuEMKHFvQ1mRXO2zp9
NU8u3odpa8/41d0bHb0yIrcHfIsjBjJoiu0nTHNU8xU4ocQqQ9ec4d4E2tzkU850m5FxjfknVZMi
t8wcuSeZ2qbAVGDLF+9bxT+TfhUuyzEEud4w9e5/qzmVEfs7AvEAKMMk9x//rTY+L6b9ENUttM9E
vIWN4QGPHbW/8p4gS1DytSqaw63Zzw6vAiwE6+QqpgC4EYbXQ6AtG8vVw58UPJ+7MUgJLlq4f6wH
NcbKWvkEjbrK0vV0rys3BVbySLkAdR1pEYHzlu+AFAYz1pJGwmtZO7cFXKgPUZ1AVmZI9PWOeQ5P
o6BVGyZenuyG3JPg1+GR3wsielSE4OGjHvsty5HOJXM0BTJK7T6X3e2O+j51JxS5QORNLl0l2L4J
AM/QoYspvviAgzbJOtc3RkoLV+LzLm0iHb427zrVbrAJXPSJo2JbXRcXr1w6tGUIv/W7WMetp/4X
DObUy0j7mT2RqRA4DawS9AUdSQEegisbMFxiJmvRajki08oqkD/tU0VHvjR7x+lxu89HnP9chTPi
bZVSzg3PqAvlJ6uKAjwFX18CHEVkyz8IRHzo6XaS69ir8mWOH8LVa4KC2YroyvROyyjqHNIpJnBt
06YfZN69n7G302gpE2zoKXmBAphesZpcA4AtIhv9v+AUka6t+XSsN1uH8bTfQILH01NAv5L9IX9h
EtSXcbsk8MW+6WVs+nr/GClrd7IAFCGM2O09qZl+Arn9pOgDTpJYppbc66ajk33DzPAGINmsZPBU
Y9QHy1nQN+jA4hMEBDmIlA9r/QgzGolMV6Zs+2Yr0Z98cdZABcoRjkO3ZGojIJMR7kKzrGYxIJwE
5WmWTGIeCXmiO0HtATsoH86l8SDYhbjLlnshaJnvxrxp4ISRLh6T0y1edfTLfOpmfg91L4E2sWxP
jPbGWGORWSJTXd76ZVKmkea2e5r4CzBJNHSPEcvu225L6mlMeZhuHAp9eOIYLYqy6lcGbos7nGXi
o4C06tKXhHWbsdeTS2MFk+EJKW49yjen5vac1F9srpqfYpMfpPmnZ3HR5mmxXgrOS5P6eaVYJVYU
XXLSyNZTnQkMo9ioVlxUWn/seZcz4DlHSkdz4ninTkHA+pTe36Ogm9b361+XrJEYEzIbnN954IQj
5o1Gi/Ngdn0zf+vOl2smLSjqKxIBou2p/wcTJ35/iIguyAM76XA23DixwP58S83Bm5kjmtge0HhL
ZrEv/2oOXd6JlxQHuwc0/TOsd/LU7iYO+XjGV2uD3KD5bW0f2hw518YE+fyiby0yfKkq+aoEYZp/
YPKWiYGPSM+Cn1daYWRtOTUWfg0w2POWyUxIZShBA/LPJLmyIndhiGYn5aSQ0OXeyhmvTmoXCB7S
Tj7oLSnvQMxU6RBmct9BwhndMwNJnxIdeRd7xjcYHbTQkXYMeTc62DKJmFU+GrF+3lew6NpPQmA3
ItgjG5beZRyXYFS30CUx0J2R0+CpovcUlTgzSx60/iy9Eu3dA1N2BrYrWk37afoqLj9GJagtORnV
J1KMgvS5vFvWdMZNiNhcYKXkhsCGaRDfaczuF2zLX5ezHw3OgBZQuCuz6R9XLfrf1Mvanv1EsWEj
upfXYxGRZkUvQ8KZVuS1lxFfgK6Vmum/RojaP2ywzl3F3qqrbM+oKJunof9HjWwlqEH/80VmXI/B
Vvhva4O8L2mpJk1AdrfoxhS53cFzW74ya/JhObHxlwSRkLAMgXPTEtNoQuaQk2uHKjdt+7dhJnOA
FLq70hBMNZ/F6XrBau/LjNJfQ4+gigoZOPFIk31KujOOND9+ITZBoSI0dA7B79d7sj9uxCd7pwva
daS0lvIN/WhKq6bUJGl+DkyA1jrvarq6iCOaH+IYcKO4yfOnmKTsMQO1Innnky9+4SGM8rT8bjzY
zDS6eW1/Y5uOZsJSqkJRAmjid13fDWXOa5I+zjH/jlTaqkL2pr0Vv+jziVLiL3xTsRCO7RthD+us
ZZX/EYUnetUgznSGSvzVFYZveZ/dzfp4niaMBfO1Lcb103QPV8vIBffDSymsraaKAPLRvvSlDTVi
2BpRRDUYCOgQCeDvP2WbMRvrzTtX+2eCBe9l5A0vEHmxyhGrtTVOvlJIlbKUpkYFBiL4GtR5LREv
7EdonAJFNc46g4EYN476hFMACJ2wFpvK0N4pkvP0ciCcxLW865t0i/Fs8CvIRWsfwP0sVyTYvzy/
KbnpJtgceq2NkT3cI8y1ujWZaGIfY/dGCWB3IGTBRLMwpod8c4qAYSmRbhWAkaCD527zVR3xkTFH
h0n/zeSx3FHuvEJIioY8g9XTGF9tfnoHv6oDCy7DkI/ih5gy8Eycz60HycaSR+I6K/8ungagOY98
tiv0QsTb85rCh2fSB6dSaWEvq0WLLBqpG+WL8Fuk72dvQFLZy8BknVrbjdwYQPCcd2JS3JlprV5o
wVH9cMjlA2Xr1sNxow1fa31IiX+FKKpkHsghLF7oCUeISXEKvOagXLfCWWo7lQxeA8MxTwDM5kD+
J6MUdhBifniKdHk7PQapvew0S7siBHGnko4PtCI9WzcyXFHfocjI4W4qb9JeeCvJc/6+8KIr5QhS
GdN9VOZE4KOQ/YlU8xyrx0m4U3jIm4hrqtg1iEshyMEgOSlcDw5SQeOtdy4e9Vcq4Re7PZIiCbg1
19wSMpbUUuh1Dt9cwYMbdQsK669W0W2omcQM3A5f+E423TaG+/TUNEUmcBgocfHdqSY12E0eUJ6y
hmA8Lkmp+KJ4kDpy4eFYn/DH15MLSOZms4JcqP49rA6JbT/68YBhP9fQXK5JNdTU23rxX13FZADl
SFcovXKSbkz54EgkUZ0gjFIT13yBBsRlJg9Ek6yy9qa8JY2roGrkCc0DXGahlA0UdOPt//mgqRDe
CkMrHBDLClwZtKDEXWVT9GmySXEAIZyM8urmUM91YAVrU6zftWCIkAl2ACJe2skGenAhjtjLNTmL
Ustk2lwNdFAvZ87BI8VdeoqCiweUR1R+eZdqCMl+3m6pyKuav1W9azaVo5p84MPJJLoXxGY1YHkG
H2ZyLZSMUDGOXvtL6DOxWYSrHYckdasWiqjPueh3xvQ5ZIQ/OsBtu9Epr7rr68GM5UTo6bA3VRMj
T8PRm5kn6FeVH6WE/6PWZCX0tErserhS2aPAMupVYMvdTb4yqrZ8sDzyIrTrB5A2chjgaKTvBbTV
ak2FRD6E3Ql5uniJLhgDE/TA7N/qzgAET0OHZ2/+NYVv4wB+1/x4ltzewPUlYm9ux4AP0STz4ztq
H9UtUQWQXRmNGYD5iuscXK35s2Qrv1O43aVoEwBLcSu6SelbeHMg9fe193Jv6c5gWWyfc2j4WMoA
dyDcJ/yOAvjMidKnPW8zjcNtyAf1HKas/fiCzPGuYHSt1PBSpVM7MxrjZxxz0c54vCvDXbq0kVuK
Nt0UurD5GfdJX1ofZtYSDQlJtBeOfJMUmS6udgtyvYAqW+BfaaYAqmafCIR4N/o85JYAq/Kq2VYR
Ja4LPb4Kwc6xWi1IAOFJR8Df2l6NTFJ2KSy830tejSKL1/ExrCp1usXKDjXzxlvkwQ+K0ozynJx1
hMpkozeGF1BNrPwejUuJgdSH6XWWRXzbDLpz4MOs7On62ftKBfcDQYSIcn+N3BEth3hgF5CcxGsp
HXDmqMAdjhgyvzTmCpGRv1VL1mV3iC9X2JYWaPv0j1TZ6VVkYwNtT8g4hDqXZKIcTDY4vTi0Yao4
KxzunKpx5W4d894CFd4Cd3IycDhNheENwC3SHtgnR3JhHOBiuZfqABfdjSoSAmsxVwvo4oZJ0eU8
WGTKEi/z9aIJ8hrm1EBKxxsPNMnUqOzmjs/+mtfmkYFdKSKprdCcwxD0A8hxatVmSVEK67/bCBq7
VZh494dsZY76vLGfPopnUs6fNqawCRX7p3hS5jFBJL7ytroXmWnu5gRECMwbn0kVb/2wJxBw9XCi
cMMZLF16JdYqYS9pySlPqUGUBhXmdRkCsqa1uxeGhe6oISSB7a2qX9oPxDHrHs6EDZO6wO5RVa7q
MtDXYWoK/d4VGmUlqb7U9Ibxf6LOXOHk628WGnBekvcniDDkwfRpy89GLwCdlhypj+jRpBgMW6xf
XEl3Tty+4a1qmK0KpeZTmVbU24wI8QpC/jn35gIrjHwqonnw3F47RzUK2Dn9AsnrOZL7ylgSdjV5
087uPXxN9YrilLeSlWCkh9jIOeRIWX5uS3eap2tnlyqtaNc962mh9e9Q3/jf1QQowt7Gpvpcefx8
8p4Y/kxotuH2prVjDKZ0fLhVTuMxieM87F94iGZnPEDtmvfeJBTW4s4LMYxihfVtz7yewK5yG0wk
hcDqhPT7du+SGCvLY+0hBKsgW/00YDCHmxpn0wVth+64VGNwYh/w2LVPGVmVU0SOY56aYwpeKJZb
xqN1OdbJ10KCJfdiX81PXSJ3LHzKuS7WfNk3NMt5i2TdzY1CsnY8HEKQlqs7uwGtK9newVsXI/+c
9zeQAIGWNiJU3Z6GKxSecl7Tbie3KiOS+K7/LrZekY0lBJ2FiokLSCkWixKS+eJhsX1GAVlNxX0x
zr1x/EVYnitYM1obK2F7ERNS/npCXbHsu56pVKvgrZBoGl0+siRyhLUSAi5rFjygs5TJRZzF3mtx
sfPo36Lu6lI0Cqq+bv4rYooIqAnUhcan3SKb4uvuBf5xwOV6aOBhqZYuftje/Pk5VGHdqLer4Ytg
PxlVPPlR2IOSRp5Oyecmus7dY2x2sxqaMvlG2oaQ3ToIXCytNJ8G6N6OIg1R0mZELRqImzijBbZR
imVDwyZYOqaCT3874s2UqZfkgDoV3RfWu/S2e9VKHnPFQ9fkZzD15gSzV9dPcK9ybteUv40h5Rms
TwibA75eRNEfQqQPhB77UL4rl1XqYQXV7ot4dGKJ7bA5M8hvQAtM4q3uvahc3iV8v9wEm4L7r8uq
Gl/H1ElQwINsRfTYTGktxOxbvH0iMwTUdylUdaw+7LKCbDHIB6C9aOGV8OvxK/UKvIX+iMWfBD7K
pLRcjNJhEsGv9+pRO1pcSQLU9r9LxHppMMTNqCum1miBpIwouv1xwq4pViKHpxihRLQUmD+HqtBP
TVrwx51g9KPo9tuJ8h6xpbQuCaQ7gdP/Tep+ssPH6mNDRsSSfIobAAZNb8AsQcaRbQGfWpR5gNxY
IFrg7uNxkooyeDZrTtsZzUT1017zxceksXvWar52Hb9feKkHPu6/ROwldemcrDYsKzPKwv3WrSGT
VvwVpGIRU01qAwhxF5k/PEWkFE7SNwHk+ztbh6FdjjhAbT4aJwoRfYI+MVRKuVnlUtQARnJ4l6GA
ZuB9YWUMmIZnV7tkTTXtRqLj/+rTZ9AYeJZUJB28tpaZ3rE4PXmWXCrkbaoeUOaFUBdvsHYhCGoy
ViknK/AxplZdy9/MPwFTp/bJiilKm1Iim5fK3xuu89VIJCkZGHhZHti5dZHqqqmEQw2WEeqvwNhM
8uuoUWppOSF5nkY6P8TqD/Qb+Auf/B+BfVURK1Ue/+rrfQBdTeXCnSxlcuCcLAUP3gogiTWsgJ8l
6L8ogOJ7OsLyX1CQpSkIaHqpciGgEIkLruIsK3KcnS2ySHB1afvxBpoD681B06JqU6SZOd8jiCXI
uzK5k8hmG8GZwMw4rse8o4R/k4c2dFWs/KqsSQ8B77selnKpgTScQ57QeUTT/oqbh41gWTn1BtDx
zsEHNXkUCqBbzo0/G4qnaFxPRyCmgqq6isNhJSN5U5h7AkJJYtvTrTAC4IuqMK2H4VEWmCkESL1H
sQKBS7wHeq2qldnt1N/3Udqsvb/fqyoydSRT/v+mnMyAzAMyWgeUKf/EnIEUuZ71zw+kvP/+s+ln
bU1siizvclk8TrWVUrKKGt1niU7DgoGUCDADnBU546TvmD5qMOvG1LzEw8bPhZ/zPfBtghUwFcEU
ios/u1JaZ+xW8yIF+PDyvm8PHr7DLLQvw5HDweHGDUCZwj+sxFCSDhGAzeApNfGsfwxcWzJsaXa6
FI8IfqIJguJ8F6YLgP8o8O717JAi2C8WKr9cFMCH9XmOMWe95+JobAsU44k0/mLJfFYTMJehVDkN
QHqh8xUixc92fnu0rJC0KuaSggRk4RJVlPpvNRfVQRE3E9OGCndL92hTXlmuqttQU5beltWbVtpD
Kc0dgUVQ0PsOrlzm8UN/brfCDl69bxsJuj4Z2XqaIHz5/L5kCQi2hirkRQ7Tfmkw52zWgu8n6gKG
+nqW4Zyo1NjVCx/NQ9g3DN1b5Amj90YbOICzyoPp6odi3Fbr8XFWxCVd9qzt5aIO0aNaxxjbiKwM
yU8mJFrQBOhiwjwN2w88GlsMG80OZeOBy6Nbg1K8F/hWqq1ct0gSvVBa5nyzvwqgeV8xIwopy0Zp
hg/i+knRtnJYx08cqnHpOOWxDrMvO7w3pOCnhxAnjqPLo3fukTGPU/AA6GAK8Q/ojfAEWDNvN3FC
Jc8Bqg8JGplil9kJXH6rT7uQ5q5/Z47AaHLsjaU8jbnO5KS60IsWQ3A3g4t7+8amy9bxhwWmXj1T
8FMJgI4PTgTGy6uRMJXiKLCvByT3Krk2cmmwY8FCua7a667kZPNs3xtOKM3UO+UpwduSdIntU1EZ
MxOfcQ3FNCCNIMeY8gonzInI6riPeUT+vIbLOGYK5Tp0y+rAdCcKXGTfmHca+sZSDqRNv3Wn84/f
55EBuICUl1AXddTXGvKhy9T9ekYQkn3nVPPB24NluxTTRoyVVM1ISV6kItfYE+Lk0ERaV0OR4cZV
MvKQiSvdIEe8wrhjbYWvl86Xc4cxiCWbORZep3BPxPwiZd6fQFhm4Y9UZQIZVKgD1rrLTJMGfbsD
VTsBMbuE6j4BZ6vH1hQrWyLeVW5P9wyOqPFIP3x06zn6Edl4dypzhMbpdrPaSg/CA0Iyv/fGlpuh
35F4tv0TeEABr0iCYxFUL/l+EQUvf1NMsXfQgmgQrL7PVZT4IUzdRHgRb+/yvQC+TD9e5NV/Rw6s
oiH7wVYNxJ58QEhL+2iLYOuUID3X9ZyIcv5DaYoiyQeBVRvCMS6Vd5as28uIoMj9DgmPFJ0EjBNC
jXDw5TDLfalSR3FdubXaLuEPsmM/Pp++Ea7sKccrl3hqGKbquCKL2gdZXyr2tnNTmZR7AkfUxl+e
wIfau575foeilsfSi2fR8OvVBw3TEPiPLTUERAm7HY2+Ry8dEDzfN4JUd7vWPn5dUfvJ+iiGB7UJ
cOTVZBmRsewayJSQZ7nxnSP1bMxol6snGH0l1VviaI4FybTGSewW6zkTIwzGLj1OgqD+i/CdBp7K
GkxmfWs8D+gC8woVHfaH61ISmCFZHbfg9bcn7nHqb4c9ZDc0sua6pnCcetfGi2hOLNLfHvjBnGaf
QoWp2rkPFKXo3MVSriv4H3yJ7lhnLvunV+pDf5ocTh9ry9NHwCk1evQ6IDD14wmzDRTo262c/Rk9
Oan0voyPIxdf3XqrGHKDWpmWUdgwg+C5ybaErhVfxj/WSY/m8+mMpNoMj9Jd6rhxvaBZzL0VhFD0
fi6RFhBxoJqPu06ONso50k7yZ9AMaHWLH3QBpoTG+lB3E4bPVYI+qLYEPGK4w2eWV+r7pVlCFQ4u
mE3l/HG3cLL9GqMKfEZtdM16q+/D48ggi2j8qSl05k256PF4WU+A998vT3xDxXrwp9eGNrNpKEck
w3wTIjgdtaDrMQ1LvuVyPsE/EA0mXY1g6p9Ynzbnu+vsRYDEfdKtTcuK9IvZKA9+2KOHF+B5j8Oe
wpghifRZgmhjFrG2nbVvc9CAT5QW7g6wrYmipqCv3TAPyTxJ8Fk8WaKE9hauvYRsnP6gyKev9E7+
OQYV0rOuWzu5XwzUSe2UCq2aVVSicJ5tEpc2DaIYWGqvnrecRiWdeAYI6Z0ULXyYVAuo5826bSFF
1/TP9LYnqX8WwhpYINf875K9uxxxRLidY3DZHEEdG7WmNcRusO3Tjzwgmu4xotaW0n1dE3SOWv6L
Xmx6v0Az2K5pQgko47y01wDQnbYQ97nyX69AJagf1+Yn0z1nihlxcWTkEdMPU09Red5pXPiZfvl9
Xiv29aVDZ6OlXILdTQiRPWPC9v7/uThVq/u5Hj5S8CkxtSRHJ6vUjoOyPyWswdoGBAYFeYOT21+K
dN3/pZEM5VYcWb6nOdvCH2xy0VYp8f+suTlsthUutC/94zQNg92ox8JWvAvb/rt1djeHfmhLIyUr
UE/tKE4x8Ejb0jCsplRjO+W04lRdnh1DhoPYsFGmYRfzQ7dtbOV10lWl01QoGcQfDSUR84N/2xeD
0bb8OIX9lylZnGVDphIdWNR88hbg5AWSc/1Wj6/xyyduJZeoK1CKa6kE3nlFxZr2oF4CB0PwtYai
vWjVg2As1Oyk0sfoOPQkbHcEOCV15VOS1XYC+KVfVNefttCoglbeHmHHhrg8aIdXBj2E/r5H1E0w
yp4ljufyT/63E+q3ViqiN3axsFBTaYK65t63fjIwpftdRSMpteZ7Qm6PkSR0hCqBL9CRVOyMhGrh
a7NSrZMYl5n5yV/V/mLTooNTfOjuUUyRJQSQfJqCgq/d6cRBOTULC46KCGGbsSXLV395K7Hgi2Jz
ULZyYZPQDSTFBGtIMDG7FXpujX8x+mlGt6UV5Is3rkP0fFN5DP2yZPg6Tw8B9lxzki0ap46EeGlh
le4sL3YF5oiUN8Q54L+EOt/mRE+4+2EgxvWktESJ3SvpGRDRogInwra0MFFtwcdcNbKC0e/5dt6X
aco3Pnm/HGymtbRoiQR3cenagk5CbzrM+5JF/Ehke5qkebdv/WEwIBJxMgDytW1QHGhDy0qwIogC
FgkMPH04+EnyY9CimdJWuxsQ0I+EX8uXaWPuqOtJG0NbEXwP1WUKsKsUCqE4bvpGVWxAQGsUwTdp
9mutlFymO5CwFyaw+byPvvgr4iUbmMwn60Z4IsRNUDJet/lVGJlI3pwIaywHNzsxefJWEvIP7y4c
Z9KzO89yA+8GU7buDdCdTthJqGKXmhbTjaBsc/Z/Yau+J2W3zRvpYzvvlZhv/whIk/TjmdjiWjEO
9iwTjIKT8CeOAKJPpwxTVndtLHUQg8nCuc1BE4wYAqRGU2mz0cTVLDswR9ltrDvO9iQyy++EgCeR
DMORkx2OHwTpjOifxBp/DGgqULG7R9zofiTZULnDtC1ZmExoP7AsdUmnFckpXk4Vzs86B5ipWdlP
Ix4bEjsMZd0aetnKODUWaMlDlbvAc3pXJ3N/+rKtcsETVUV717LrTYYMUFWyQgRm0FS19hMqU6hy
K+H5z4ECvHcczI5TspQKneBXYKOKeBOwo+roNW8IoubNDYKoHqj879/r9urSFFqMITbKPFrVDM84
Z5XdIo5NPbWS+N1+CTMWCaTU01ssP20rnmlReTifZOSh+ESoYSli+KXlooSfFi3O1FT6UMM24vKE
tv2La/0DHaH+3G0FncLvCC1Hy9NvU/pPWGzmseR2P2FIexZpe/CrniIsymjEatn195V+CaXMl0fn
d+ti4GPwkqkSNofOS7EKuhJARpshyOvXxQn80BZD74i+b8n68xHR3o1SgFunUET4rUL3sMktONbB
Niu5IwF2EFH3qEXyG05Jnq+yCtXdRoyWB7Hy3UoROUcu9lwSzN5PW3QjzHjPzUrvQPwM4mpVtNjd
5ydy2dZYSxnMi0SviekJAWLNR+sD7OEUC22LIaMj3tQK7lAZZPf6yJqdsZZDie8W6uLR3rU2Hbb4
8Zj/t5Yz0kHc6Pvc5bWD6RUmf/rXqTTDGlyf0+Z4b3hfArd8oW1BpKKJ0iQzIM+/WYWLvTm9wkez
HK/tVSOykh+DyiwpjisxQa8g6/ztAyJG6MVvhGabukZWrrYyae0eI/E8G/SxqTCZtV2KTbY7IH2l
z7gSlqLN2lyZLI6I/BwS2pcpeukWsM0bYMhUBPWNLl3c54GNvrvIX5AHuE9pSiOeQVt0N65Y44k3
gY+BGGSZQx4/84NQaPPZbr4gsRlRdDQE3VyFjCdtpL9hR1Df1uBMibdtmCzEilkSVhJNIpShCFko
b+0fDJASI26aiVr/sDXsaf3LnMX4t6okVG+TNKFJhtOy1xFMEUYVSaYa06W345fne/16UavgQAav
QAmuwIu/IUhpK9XSaVT+h9z0zT03+FhuV80DUqpwYRVt6pWa4eMjGkfwTOcl7bUbMlPsrcMxKBAw
iEUqqhR2d0uVI0oX0rjvUQ03wjnjn7dZOD5zd3oFX2Axo3wvxZELWUTeMX+qgML7aQFxP7Qs3dDs
xhqfhzTSucvQ1d782EBel0TyIdbfidsZb22pMI3xTQH0SZVUWiCrlUuGsnoXLBWVr/nDsEh5vRAY
iifOAuiZP8CPsJ9BVQ0kLY53MZd+77TDbfGXD31wE1AxPgs7WaOn/6T+LiN3kR60Er4CObywuJTA
vbxOjMvy/bNMonv4jVnETD5aJ4Qzyd5yuvMj+HQD44syoBwgEy+9iyv259w1kSLqZKV7AKI0F0gC
Zg80cCyOkq/wUQobqh8J5BrOjhwYOfoIF/YWd5YXsNVSFVf81Lo1K3ASlfj3j/ylS5VJJqnsBCuN
Fvep7+YRxYMkmON4PfcWcBzKXk8oG72e42zWK4RdXoiLVpTkoGUaid/IV0WoeigQ5tRRDpqmhqOF
l/5cGd+J4P+m063lLrDF1UzAi4A+F+u4Wvf9/DHTjk1hfATujARGKXw20w6X/nSWC5t9x8+fRrFU
ez47qGDW8KdQVd91E2OPYmTSLTs1QiORvC+tpOw9L0CQaujxq2BbwnoBfe6PfyRpkVmY9QjtHn9y
ux0qX0AzfRttoc4ZMhnp55jHTwwyoMZtZA72SpPbkoRF7s+0p29nUw3U7x202EHNiUXrSZHSr3JK
+7ZlX6MjwCGT+O9bytEP8APZEHBC6hJLobX8NvIWaPeusDBICSIXVniCxCbSsFTyZ/dbsJbDcSCB
02mNMWCpgUa+6ikeL5rz93anUmR+uecOPtRKLw/OwVvg4ajuW2jvC9qibDKVxNL4q1mXuiryIo9k
pETzjsxqHkzIokDZGVcr9IJTh4+ycMnAVM3YB5zb52RFzXHIYOvWlr4Lfa6VdYLmTi7mb9RgkJMF
tt10ZiTIFrXbTCWLc93xQexkOHJQjFkO+mneFjT93vj4DHdIpxi2iqTg6xqy8speicOXcOd1ixol
C7yafaZ+fC8IqfbhQ+XkQ6PCIE3STatubbYwyjFGEOXxb8VqOvXiZkP8G0up9ibYXE8i8fCv+AD9
UQ0PGMYbEsrC8vAEBgPRzdD/QxaV3uiQeoc0lE7F70s3nqrT9/TIUUeWk/Tc18iWrN8Q8sB70RHy
i3hj6yrufgegE+p9PKVBfZXrJf5jl0OAsJGwlRvF2iDTa6ZYJYylqACWH9wqJd1VI/JtGaKIzpWL
XPMzJsZzITKk2/JviAXtCBs2p95tZ/7JQFGKS7nVsxDpOCbKUzoXcGPNttSE56ynUzSiQl4B+Hvm
9C1+gNcmyJiO06EA3vMgIQO2fX9T8azYxdawF3wLtda+b+RAeQv4s60Fz7amxN/DDwjRx6PMW1nq
E+nysjQDR7gpx3v27DAj6mc2hAbgFkhIstOEJ3Kt3mh5jqsbW32aTkaJgQsAZvD8e5JAtbM00lsk
0x2c/pAWMB0K5IH7sdv5P4k6OzpqVfodK+XAp6e6vqSJnHJ0weJmBYuxVuOO/1yM4u876jN1P6rC
GzkNJ5A45Z1I/2ppLLrqu/gF0ycWl1NjQYX39Ewvh61Tyt/le5VZlD1rtTxyyIPqydicgzESfqL+
FNnyftxJUyLz0y41RhsbvIFAYWBd1sAl20WJu4MliLZvKrDnM8c0R5RUP5eF+zsWZdttMDEb3Wd0
g+J9dZm9qh9XWMbzbz0/1/TtPnsC8EkKNzVH//sjrg/bEUP33ioVXhSQLWh1stjFPiqLcLreBlBa
6TYOHsjZANc9f7tx4DpZww6PSr59OX2ZyThyW5KEdhnK4jJZ5NDyvRDEcLGdmEfyRUSQs2lWzDXB
HLWramoGauMX6PYjvq+g7FsyzG3f/fE7Wd/W/kU0sga3pVPvui+5/SsH82h7tweKth7uf6kI8pEu
9u9s/gKZJSjLhmpHB7mNCEvuEAsQPlDScUd/hFl1+3eYZfh6jrFbqB2YkrxRbIf0rz4jgHI3Axwi
JSiHoOfzLWRz678s+0U3j7KvT+vbW776dKyenvWrw+ELmO+rpYncEZwLCcqa7G18sRGF4ej32qc0
wOtwCkxUIKW3iE3b2A5lgDxJjnvTRBwdu6nJwXJQxyGprfblCVxDhkwb5rDMPUkmKX+Xw0PwUVLp
eo1fiH2s1szMKueA4hj4YOdvnzZ7mMI8NmmNQ/Fm/jqun4YrSgzMgv/88kawtF4kftC+h1ySsWTO
GbKadGgOAcMaMmaLAoea9k96N5n9EJiUodhbt5NlNJLTViGBVeRmbr0HXHOZeHvhR2laZMU9wQUl
zLtnUnC1CYtI1cX3k0TDIeBlBj2xfzI3xR7y/8VRcBYQ7OwnHTpSKtH7+7Y8fqFMXhzaDuOSARic
R2MzGERdv1MkXgxsE3YKWjgZxwkJsHdMXvYQuar78R/rOQyidd09axWTSy0InLOZ+J2oVvODyasy
HOMvBvnsKYoI6d5zEk96Lh/lUb43UIf49AJb+xufgIZKKI7HA5sDxX2hUug5QXKZ3kjkhSaOJRGW
TEhHMOWOekNp5d6vKeVU+GPO/2Q+2bQCKFFZ2a4rjRXrnMIKNex+FJ+hovWqUfbPIm2rdJveKMp1
a7PeGpI9Bjmz76oDikWMGdieELgHdiOoJnX1guJQiHO6p4zU1QxhlnTKa3+ApZQ51t+eet/frhX5
GVTv05DB632XApjvWlQDTbWJWzM46DSIGvTJ9yIDqKWL3Ur/4BVMSzgvnw4myODYF2n3nplhvBFm
qw53rw4enkrTTfRjYTUcRKcFeOdpg6EwstK+apHDefDpm4S2BSgHVFDGEsvOLDcsV1VjTcX3zyJr
siMZ65mnh1MDvDVzAQDFasZEGgsIwT6BM0oL5E9zZrDp9ssSYvHLXAiIcr3kZw7KxD6GrYZJAAnT
m7U3A8lzrAPwZwGbDEPnnhmRyS0sR7MNIvQwX+M1EN1oYqJrX7Jp7Esowo9sJjA/worQtw6RyQZ8
lkcKTvhvpV3YfNmqhZZt5wQjXQoV/SWpQ2RJLHeL0RVNbi8vR+wXyNXykCl39oJT9JiiODOj7XWI
Z/qQhdpSsmxtL5bzgJfG4IUUk0JbtLAnh89pJzTjvCnYHZxLMOWeGTaUQPRYSSu+9rEfVmquVies
XyxJSrPkFNSnioWLBJ7o5xZKHhqLbJov/h0HX3IHW/6bXZIsNWZmM9zq3hmEgoIbRlEoGqHGb2Rq
iptMBt9keKnuFDJrFGZoCNDRckjx0uUWCqifKM3POccGyPz3FMjSew3oaUdQJMgTaLVFc9vTTkxy
lttR14+kguM5RbRmbctyva3Kfumi1iDewq6tjLqC9aS3jHgCQW6YZbV/Hq5glgV9lzV85L69e+NS
QLhU+843DfXoVyWrId80hBk73WzkibdSJBqzyV+LQIxhIVQRH9MxCxsE1svW8iVuyAqJkRgB8oxl
20O/WJ/62P/y4DuyBrimR1mXMMHHFklxlPUoNf8zBDSBjIhsBYZ+799gTCbF8rD8lvxNbm/GLZc5
TW1MlowA+H2ZkAfuVD8RGyz3LdYBfF/jaUhwkCh8waEtomMM2iO2NF+OSEbj934JfSUMwa9RxUmL
fpdaI7X1YUU+XJRnwh02ZqpWaAOdvyMDKHDgpZyUmmG9b8KRmADj2vXDr46cr0Ipq/HHRDSTqpEZ
/iWK39N76tOCRFLMzDRlZJ42qZ3aceoxTE5cQdi7i30CGrfkakNeEAAnKIICvO+IJzky6Jgk0bWW
awDVKp0xlSzMjaWwxNCmqkki+L6urwkMwvAGxkezAArM1spGYQDdgqLzH2IvCg7hCMRaEaKSnU/V
153q+FE5ZXepyiwgBVwLaM9D5D9klTg0R41IRF0Qqs7450NRCX3P8KjZO0lesxj6iL8aQD45cqRL
BZuGzlQSKg3/P/cRE/c3co/zlOqVDfGbvU/yklsmDCbn0tZr0ZHB54TmPJXOftmcKbUEi67gYyL7
BZcpZdDQmYdbGoE6x8RT7tLV6OXeUE/f7urfRIo52UUaDrXMqEDpxb3sAANyvJriimzCtJk1vxJZ
5cYENRYfVikzwpn9g1DzQS3Ry+QZeoT5nfn1B6wq16Khe+Ayxmx0cgE/OK9DcdkDaPJGOm9dQpVI
Zk79VPzFWxAoYSWyd19179yGdGTkoSzxfcnthCbOwc75zHP4663F7pRp3eWj+Crh8qInXGpf31F9
ix5gaZLvQOBTAroo93tyPLopEZgcP0ghz+cfB1fckgUiJbpI7KMT5FeQz614G9jBabPuxL0OQDPV
aJJwJS9k/0J2O43AMA00gqUvKCCoyysBjsumeBlQW87j5Mite26w2ldLErM9U+EQwvZTH2eMd8Y4
czGPLzjdaixiP3hpcoiq+JBmyPTcFbsHzR5FTRitOcg/RdzoSnWZk6d4kuFHJwfvTp4/AiPTMPed
jfvx3Mt2/kXahOkfy+rYqWicOQUfpA+dfE5napcR9i6Q6hYcb+L5IW5+g3OfsF4uac+qibJH8OYA
N3OYyqsQ0qeb9UOLcKgfKd6kUeptZA/8NwgTL4pL+Q7rqw3ExhAeYASr8rRZfuFoIh59KAIkTUnW
zJ5wNwktpDcLua/ttBI4dqR0XraHMQFkCF6ZJtQegub179k/Yf6XrNR0qvMezf632Qugd5MEZV6C
FwzJ6cBQpHc/5cu/Ni1QhJcenU/PQdC9DDlKeL29eKXMJLgtFRc4n+l2cazk78LA8RTsRsPLW5Bl
V+hnLWN7EdD0LvlKAUA1fuORyJ9sEVs8udsKudytNqn0rnLXPzE+9rzN/sJAd9qZdMstvtORV9dU
41PDbEA/CZ0UQDHO08p1FpvKkfMsxtIVU09XNlSKFuknJuZNigZFYO1C1ZHq9GQC9DtyvbEsYjn4
OiuaTyI424dxt6BFPZfsbfjHDa9nw0ZB/TUkqgrsdxQwOIFOzGOen/0/mNzeD/QdRv8i9nLNOrFj
7vA/4TFr1FRC+Y1qHQkNoEWa8XJFP9CX407Tg3reZ26SlUyQrz4g1NWxYJRywTQhjDG05IvHzFOM
4tZH7PI+G7QJ/aE+9iAYLyNspRueCVmrMojUwQOs1n85QIS8WFQyI/jk9rqkhY9f7f4EfW6fIQzr
WItLHSgPH82qgK5J1fOYIrHEs6SXIIA1N+7aC+vBw3ZRxLG1XphbBw7CF6Lif+Wb1oy6kmg0eYOl
ggylJ0l0Dz1lvCVd57d4AYVDG/oKjS2b0GkPwSdz3CtcJ7YsmZS+X9vV5atIXW+AOgyZh3HrrRRk
lvWNqk/U+yO9OjhmSr8ag6ufcs8imF861YQbil703VE/1usur4I7grHXMgPYJ4MdNC3HsBYbB7eJ
V6ZcPMKi3AVFl5ayZyOpPhanQnVNd9it74U7CqjnGda1iJOGxuh5w7H6Jh/a2qUTqE4VKfCqaYuB
4Zw3kRlEARwcelSyz1wcESlB2nV1/t7nWbhnZjTUXPnLe+xzbRvf5+PwKhKosW2U6BQ41I92qufZ
l7gbBYxt+HWmkA4W3o3cV5NOeS/WlT6WLknI2ibxgYAbDkHMa213LGgAaqbdPAigFOvFP+NoUwDA
XTYhpNa3Hoi8vdLCSlxP/K1tRJklR+VTXrb7vcRcDf4qrk1Kv1fDQIzjH6BnkQelRwpS4ckFCGlF
kHjcVzDpL+SqtSW49ksrOWgHNvLGwxI5gTzNAFW0qvbRkYfOAA9gpRg34an4zngGjTlyM5EnHOu2
qYUmWcZP+ju1LcOed1Iea1Mv+4RVUW530TjsBAPc2CfeBk1FP9DoA4pbHu8CeDHKS1K+ExnIO4Wa
35F4Zl2B79a72vqobSct+I5lHn3YIiUIlEn4IoxBA9YX2acZO3rDSFD0j/67x4k5CbAstWhJyw3C
38tmejWrXtj9wsOlK87l4MsOsi1o4smRjBR7Fx7JeebJ52Z7EoZrv/ZrzXNlO8YccnPe29/h8f+K
2zjKDYE7cty4mUOra701AulE3PFT07EmJ7i8iumCy69Ybepb/W6v993XfnyMhFrWxTb81QOSUOj+
9B3C9F3IEtjQpVXRuxbzqihHtA1u9lYOBLIjfyXQYYF76Le7fpsre1MJlI4ZENeMKFDW9/VejmED
61WLwlNIuG5cZ+XKWnVbGnibHvyGYe7PjNXukicQmScFIxXl/O3Z/ZnwWVeRrPZkF7sbl21LzM3N
xotrxBTs+nLWW9KekzQwUOWgF+6LVQo82ibQzIrNDKux1wy6s9Y+U5Vn/vpzT3+l6dQ972nd5IOa
UV475govoc/OSAd3oqQlPqFtcpAjpDLaHekdScHfIpMqJoDih8//Qg/BGWClcd1BGnS3OYGnDVbE
M7F7eOOaR4oLF3cBRouY24Oh5KdJgyae7ZpiiJsvPpTyD07oVTZtcBJmqVi0/JwRx9Wqoq28Gtvl
odbR6pOTWyTtjA/mEL+fbkGmI7YNJFOE2DucOwpLqgRnUJ9u/7V5WYSdKcnkPVu90MbyqPEu82yB
hPd3i3oBD44OqjBze4u8XNicCFURjI3CoLlaeXa50m5i5tmDQZ2x672KXr4N/Xt9DWLaHQCh7SUF
UtU6aQ0a96W7Mi7D1NFAuCD9a4p6ifBTnl8H6TurwQjgzzl/IzNDm2EiGJSrIGLbGeU8r4z9wEAt
kPo6bSWh5XzXJgUbd/86creOruJaGgVGvSlzNmcO3AneVuPhk7P/fLF5PEejKxsYMIgcUZB92Uvw
oUuIjo8k031HP3oSGihRDWmNdaOOmnDsVpIhkyIZPJNOXsT4lAnOSzesWfyFmH3jc0Q1oR50TkIS
NekdgIudq5e5wnii0cIX9ON7pI2kLw6y+1H9kLhT8G1wOQzHlbtfFhj+wpl2rmF4XTBvo2vrNel+
Bjil1xOMfKCuSrxo1RuWYHRxhF5h2vGVP8nnnRGjUBCm67SuH7oPKNIPLO0KpgIi28KhBG0tWjFi
zCNkvRqKfNxfBwR6hkKwpmePxP25itgofLGgaVgbMC11A2mFozOmpwvk1ykYkFhWVmYaGselOXVT
1f+M3oEegmtqYwPmF4gd0emCVdg7bFzy5Ydd8ZF2fzt5Swtk6k0raE3/7h4hECTHGjq6HZODI8vG
2j4kz76a7r1XYIMkgddkdLnRhIKSrUzEUn1MHCB+/jMFhOuHCbSS5yITtM38g14Fagjo9sDN94D7
sBF6pQoJrLCy3tPiMFdv1FIivk2Yn0kDJLX6hyO6320whWDwZv7jyk0cy5v7eFbkzdBJO+Hm3Koa
9ZT1qMlFPsc3iu0XQc2k6LuHQgP2ddyjh3JJrvUeYYxRWG5kS2g0Fn1Hu94kZ0WYTJEdtw62hujJ
zRXQ6Qb0psyrEAj25IxWqett+L+IZYoNLgch+/mgphI5yS/dnLs8M6KFimBdDoR2P9Igitd5o/mi
HfSW5zhFGzotWgzaL5A0uSDF+89U9Hr6SP+TWxDNUB22o9NR/2O7TM4mA2BGYzXDVqqo8Nfcg2fu
/lurynIG2hgKVQWIkhRlCRfFnGKKhONK3N4mmL0eIn7tKwtQYw7rJqrU697e25VfqrHioarkC4HA
rPMNK54bJap2wfouOuJ8IhsJbk16lFcxFODwI+H6rQ5bObDhpEDgnxl5C8wunHKtleQQE9WAGOIg
fE1efOGDjkqIKVb1EkTNQBm6laiU4gEi+HyIYoEucHQp/bKStriQPd6CdJ60kx0zSB/4XRRAuqQi
JoqmP6vwHDnf1lfgJh2gXq/uyBF+EZGGZl3VkpTOoWP5a+aGwG6eK2AoqM7Lahyv6UoQqlYjsIR9
bKp2uEaVuVIje8/uHHR/qQN7vv0Xc/duud43V1CWWE81FWo4rN5tBfw9hs+h+f3tpR0nczZXJNvS
9kzX3bBYviYpqFaO12yz6ISMQruq9lAcAa+unEggvsitGwgG2YjAbuxyQVX3pvLokF4gVHap5+zL
zYekiVePDHWvnmwxU14+cwZ6VFdfA/NVoUw8vXOfOjpi6kCjBtN8QCzMxu/QBaccCyJQRuJNwuMg
JD9VgeCOvktFY5pnGykddyjPY4YF8RwIaRe0ibDPdG4pGzgZ+IHt4p/UiJL1m2ZdZ8TTtiUMxhKJ
8C/Z0Rng0QzBVUvWuqdA0FvShOnQZBJnvg3BJpws1kTydEAW0UbaLYOAXpEtiHUAbOzApF3U7t+8
2WZtzUipNCKuAHv4QDxJUUSJmNSxdCHx/FWizsRM4AGgFkXghOShy1qPUxBo124i+pUIMKKFwZOd
p1nMDpWZQUY0blWqHzwA052117R7dD35IUt7xYa8AmOMheXXE/v1+4shhgP6+QJaOEAIl8GRHqrR
FvxcZ4LjoaXsa0/w1wqqpFVhrqCqs8j/e+HLJEZp6IbBiAv9OWQ4UY7EjA4/07XtLQm5iblXaBeI
YhaQximD5VTW5fc25B8HuByOZYsiT5IOFKYoU24pFun3TzzLJLKAxImV14kYuSEjT/Fu3KVFak/5
A2/KLNX5CIaqKQsJRg+4ouC9cjByGHi/EQgmfvHqwsOHddcaFDYBJlNceD7lqd/VO8nVa33TZZ4C
DYePGVNnrRtC/sCUMsh068FWDTUZDzbdd75pxTJacPATfuvmeDQwZMsnmaUGbqE8CVWWvHIaVt+H
iH0POdX3ijBG6TfHmO14B1sxvAxicRs7x+1+w5xW5gHHaBDGXEyvT/97SSNDDxJnYvR3BZ5AMtsZ
Y5h/SdjIBxLc/WkCUdITvkFmS7ZJ5Pg4wEDl9QVQvN/XKRtNv/29wTrHQ/NcFPQGJXDtDuJq5hWJ
Vr5I6851v/J9ux+5XShhO5Z9pudqvnkorUpmHDvUpu0G9kXCkD+3WBUgIUwA5HN7gl1MKN6vP5nM
L8TT5UZmTEwmsKgAIn3/UBzoO6DRx/cMvT7PhFm85BaYPKDvpWWFfJVWPrbvhr5Ho+khk+R+TXsX
1rDhdye7NM4EAzhQ79fD7x5L+bP6hBU37x2vD9q8JxIUxxcJSRriScZRGe3dUFoeKEDdkdYiVq5X
UB4U7vK/4fLQ+ueWDKLu8OpqpFaumWl/VU68RfOgKKW/BrnJkh0QnDmv5Ss6u3SiFrpMk3swvkxh
UZ7KK25AaRKjQK/NwjR07Nypo1HUpFvLr6q56/t7MDPPf3oHqoKROwJchOBLskOegHkSGstnNv/O
pE2Ru1rc7w74w5MFJPIYHT1a5lQmjTinsVxxYu/jDGzq+eEWbvBaGFUnATgjbnC1nXfW/aShvVkZ
+h7aI6HPE3ZJM7natDeHBmHFsZlWSBoYAJlFhx/M1L8ZFc58e2na2F+eJSa/KI7CBQJtK8tyzOY3
RA7/x790LyorG1iudIEkRBN9fptNCgHlKZ5NE5/CdQrr37aU8z0IJB1CYORoQgmTB3ebmwI8PUHb
+7M6EBIHYf4dFNR9n2piy2InmOAVupsltohbRkPApFNT3eV0zJqPiZbAta4wVM8pYgH1cp6jkk7h
jO8JMtXX62rmZ97jRhh9Z6OMh3sT4fFIGLyGIX+/X0aCoz8RPUyFYZdXxQACiGHO+NzUTBeyD5yk
mrrA3ktsttmZTtxQFhcFzjFN+Mmc1P0AExQDfHxFExhrMkEqoKywE7RFHBaUt1tpvOCQ7QQiBCSp
1l5jT6au7f9jUmfVyIb/UD6VRCDadhaUtNcPhdtIcX3RW2ijMGXRdN2bi/ENxXCNMdcY0VKbsYzH
NEEBGdLK1xHnyKRzdX+pYewW/LgKu3GWL8RXF5iX1buPxnr7wT3qvl9uTxiLDuEAAkcapbVtwIP3
xO0EKXt6utlYiPKmHvzFCe78ze9o/8ATBtTT3WdbOrUk7g/u2FWQHZTUYt1ZscejLeNeCCkS56kz
VcUdt8yU+7c3y2zU8IQUUCjU1TP00RPrrb11ovHKtjZ3t019QZ26Nwgx2o4gsrmPTyJTYR1hDtgi
yIa1KGbNMZ2llRimgrLQhjDqG0DMq/ZnHUnNm8Sc96skWp48HL0oqOS+NcjsvvnyRJHi8vzlJ2ff
lokBTiyotW4cErI/BZmS4zWcmJMIOzJ3X3IdH2qeIYBo8p75Q0pWo0tPg/Nou6f2LcpwzxGGg8Nb
khZ8fYbmGyP2ovv6s3W88q8gnoaiKNyiD+oIWogJDp6mm+kOWPQGRT1ji3/ZA7tm3XDmZIEfUH0M
ELvTIrDNi/DpElZiCjeY4OK3Ethp9qh8Pg//eze5KXLyFcTCIdoOcWtnW73ptTg6OGp/4EKMx9Bk
7b7WXgFp1usNHUR/aeaX/zv/LW6w0Tw8FGdwAaabZzzUUZ6VoH8O14IZGELMS5qWn9x47dvfnc7m
VWRxwfhJF80qis3dgnCKZjhmGiBADedckes8UBL51jBZmGZJEwTMoI1lATEDZQBaYS0SLcYL5yz1
2PVRcr3YWwbq4Kyn9aOsMLdkRHOSvyYyRefQzgsC2LuiMgsci6n2WkV1w0Fbqp7NB2BeXezHQiFt
Saxy+J506iRTOJARunWBNhUQz1MebjDIwlqxfuDfS8g3T2CGtzBAGyALX23r5SsjVWXdHdlO5d9C
IUW+GXiOvWmVU3Rp0JrpivhqNPwcNCIKSZowi9trnpRJ4c5zDRAYzibuqfMoni7ilgkLDKCKLl6o
9JpgjrhpBCcriNpbjrRwbxaCCevLtH3NIYrvEPJ1XRNMvysRGfh33WVheWaZ4fTLDlI8T1BvshBX
rkYjklGG3HsLZaH2HG+XVgO0FnUMF1jgtKPq8q4+jIJziXqjdafDITszhHR6Wi8jA4eKyozzY2LO
rDPI+nVoJnB/sXa/m/Q9FqbJbdX6rLN4lJq6xeUqRZneqNTShF7JHF6uGj7C7YMpbDubpjA3l2a7
YOmJ1OB7CI80CrPWg0YpXyb3OfGmm0uvBQI9Y2VxwoNmgSCE7AnX2M7gmxQS90zpDrnv1BMNQs7V
jt7FVWROxedHH4itx832ro3lBJuh8tJwX6/JasoFmjg1P+9072NCMjjp64Wc6SCTlSODE9bAwz7O
S7QzfpqedZvSCE7+6Ml1UoJpEMP4JN8ZCGAuoFGNNd7OsY9NNB6ZEBRL6Ixia1XOyghl8RSZvtgc
I+pxKVorRsCl3tU51zw7rFuM+wQHvMnp8UUtEZa99pksjp0Aa7EcRlnZy9fSCeo/yZ6CAfxZX3WV
oqKONetAQGnb9UYv1lx6YREPtko17/B65IxCpyD0biOlDrvU4jLEJ0S/zdInXLrqc+SFCAP9GvzF
zZ2r/ilVlLd/89z88pvYZeSBCZ4UCiRdieq7LQhCeDKRC4yUH087C58U6REzkk2HLc8NDC3QDN1p
bKcF+mdoPq6IhrPwnM79JgT1bPBGpfdQylTIagDzf0Qqvm1CE8Doiy2hrvyu2C2ZoULrUmSlOS8A
Bh3+0bDVpQsIn1UD2QamnuAnYgX0UWnZ4oOsOG/JoTYE1F9u06sUh7jMqfR9q2Dfl/3778INKv6P
qP8xQzQsYgSSrjAtVrI4VcU1P01XWdMnak7ZQgK1g2rO99LyILB68TzyK95L5kPdbtszLtUbVhUu
XJskA6u2mKzM84eX9JIFI2O1S0DmJAb5HywB1nZy4mNEM+iQ9z05KZmG0coo0HSeiBDBsSFN/Pyh
GbC36Zh3eJUk59U4NvQbaX/PKDtIySpZzYe87s9adSykbHFwUkx7MM82QMfakNHT0kqQSFfl9Ebl
qov0LQlS6h4z6Kty9zzzfFQQTrfaoR0qnZvGkz5x98ceM0PQh5x53sA5kYwXpttSNM1HN6DB3dEX
BMnsHv3bBmt75FqUZXzyVXTtMM/JMhYsiPyEPoEwvzKakxSQqKVwoiDtEx0CDqqG0SdzS2HxSAAU
q2DyRtckYEMbX78egvsMwoFt4cv1AEGQ6RuPu3S4d9vJINuT429L46ySVCsnzriSUUS+L319eOkt
urD0H0ax4D1IBTpk3M0BjdR93PrmOELeCy43kzhE6oiVDqhePCTmblKetI29jx49FZku0885V3pj
Vk5XSHQAG4RatIysckIjVuVJ3VVqmkAPiaNIIHgFVXw5csCtjijg3XC2X88WEkJ9Yq7F1Nc4yM0N
mmm/+BkaEr+bPrq8vqEw9sw/AB5YIcYCrACe5BCFVvO2g2B2W6itZkPIr+MkIEyWhaECsQ/7+Iy9
6ZUqpzVcwVpdna2n1Ksivj1BkEBZyiGJz1gN2wY67zvo7KBd3DAOEqrASSo0qgfdhaB+CJQgsUJb
SgA5BpTqK2hx2IVd57/XWhgyANmECdWdArPLWAPBYRcBxAAc4M4je5dbnytTfdYdT58s6xNObwYd
IaAPJUMS1Kmx4j7Td1aoZl9C6hRo92CuLqsZETWM9iRxWl8t5H762MgnYrBc/fIG3KDHDnlm0ZlG
QSDni+xDtddIN6H2FeCAoSjJKRYiH+FlNGxh7PXROKTQ1ZSxZVZqsZ0xdkzSjzmFlvGkjv0HWot9
j86lo7wuOFL5IFYkB0QA8QiatuiHw5JtE6UMvTlfi5Vopg+g7wRFxFIDrkYtD6D8bx31kvCHY70+
rHDftSz7HZiHCQ8B+k22vtqLUOFd1NyWJgKmDVCeQ+mr0L4krLEXxEWulESGcc3KdQCgegbH4g7x
iHrAJhZA16ADlhZAAqUoQWrxaiSo0ynOGlz8jPTA2G4oxkWajuMr+gfdUDj/PJuJjX+6BJi2lRtw
88F9uHU+SfDBkeueeBfOtm+lt61VGqLiQsKuUveavBbkO9OByRdcY26oiEkYgvBOSCQib3RN/2JK
7uZpGQ5KbOhScl6hX3/6zJ+KiLvijurwyLYZdb9ZyouMeGQSvdmvt6ctU0NiE5iMV7e6qLHQoZrB
iMMjbJpGgXbeOm67RzIKNGg3Zy59Iq64EQdZm9MjFO5hdFYaKQnwIIr4gOxfjO+GLXM6hOikeDTa
O9zamh2ZnFZ4QybMWDSspKqorOKHQKyXwc/kzwai+GZD4aJcMskq9KhlTKllUho/k4NeFA0iuSJ8
udNRGSTNpRfDtxVLcGKBNGAetf392VlipGEtJC9c9Wt5aVMdTfyx7F6sej39v/Xzxc5GJ3pOEKoY
l+Iz+7vwHVnD6QjP/1kXgy6iwaIk+jTgIb3XwXdNwnhule28l/nsiqXXkz2jRWlzS0GW5ZeOj40f
tyJu5zrBz32adic9gl7prbneQ+o4MwoVrQ4o5L9G/GM4Lx59WbQ3epGalGYiLg4oh2U4KsV0TOZW
U4LIG9AXlImEtiSWsey7V+UkfF5vD7uPF8qHC4hdb8tv2mybDW2t70ldETPRr2ts1yNpHd+Icwxm
CX+Ssu6D9HmnQJLV71ZGJ5C0wz3LpmshqEyRv2mJdQhf0wSsQgMd21xlM79WpwbetwBBF4haL5uv
eHWhy6OktZoSAMda09YxAvNZZJcidHUcDdi+IXqndYW+GFbg9vkZk0mpVbpsylNHliHdrx+QUjEf
4dN0ch8CPXNersn9gxVtrIlO7dX8Amc8JkRR8hVaqIL42Oy8rAyuCUI2+1yJwB9tVxaPB0Q5NaVh
ujmxDMgJX6+KFx1+UC34MSDTgx2FGAsqw1Dys/VwtI2YBm6LkWna6CvXRXA2GfofdX41TOkiI1qa
p7dmM23zryLp1zSsTB9K+QzmTM1lm+/j5kP311cQrgE6p8RJ2wFcuDK3JP8f369HEA1EcwnXqqWn
cay7io8yrGO9M2mtGFElZ+vSENKS30+ZnUtA4MUE+ZAYQIDxy1Vjxv+gyhTCtGgGXhTqvt2TjpRF
eC0vRirRlBIOHOHtOdx/mnku+iSeKAWT4QsQeQ6zsEQrDcpUDock9j67u0nj6l4uWP54WxT5nuLr
9Wy4Otlm+IlPFgoLigmDHKZYDJFdPZOZjW+0CtqopHgnIJC9P2saPOvs29ZR12+GiZkTDx5Iiv/J
Jt2mitHEi9iMZBs+l4ohBaeUxsMrId1RJfVbIhXbhMOYNhQd52eRbjDSXG5sOZi0pBtOoBBfv2ad
ZE6Rd6+8qm3BHORSmoMLlkpKIuXV3uRznYKnYnvhDmJK86wGyaXkBH6RXb+Lc5aAy0xH4V9NBoXu
6fAX8HCumL2xeQYGIaePgaTQZIT2w9KC3D0Nwbv+tazVSxthH5aZnzRXW/Pp+ubXKLXTFwH+J+II
/PRLmu701XTXS1yNx/dRD+FEMfv7wVOe0UDTXU7Ee2CJlp9P1xNZHXhJ0mU0pPRt6uOe9jbf7OsE
4Dv6i5K4Ru3Ii3M5pvjrzos40WVJfKGe/9U5jFyZqxSfG9mDlh0vz1j8O+Z83L68rVdA9+LajkeC
8bOEGcnnaySz2O0bmKxXyC+FswqyGnG8Cs0vL6nuGBmJf6JOqAO2Udwhuem5O4KBZg0BdYKjf8NB
RH+YpR2244EQBB4u3DSYYE5/iTNtdJcCEQdZC8DqUa1VTni8JaI/aLtKqm1utVownbTwfI2GPaFQ
H73D3B+WN12IUfwGp21WfLf6THSBDwWsikF25GLVxTiqy6XKU3BsIbehj12LZD1Dn2z7pvG8Y90Z
81BLssyLJt7yVNzo0FrWIR5wJbFCQijI/o8ZzJ729GV30sQcOhZdv+F2SXqg3D/uyTfI4QMwl4oJ
KSBM+W4qVDndQeXB5uxaCJsuF0QGSfmrhuv+RoUWYOjf/XRnuHpwBqJSkqUBbBcRACj5TpCB+Q48
pTU82o677wFCVsj2bMFy0J3e7UpO7r8JdruQ+Eq6nRW/JrI11S/3J3jbQXnD5Hco2qEDYChQUIvU
UjGlrd4nl0ZAzU/e4FjeXfAmkp+r9GJskshAbN3wSLABsA6mnxTRrYHOwWZen8m/0SH7t8VCkhom
AIw04ntLvQMKCAgGBxMbk9oSzY3F16NrjR9ME3GpIjMGT1cQxz8sk8tKmj+stpJYpPjcuJ4Qv7QI
NqOWaKjHQ3cVM3iWsslFUkwTFdUUfIPsrF6268cdIWXUAOXIY6pwahqIpQOS1+MqZ2dxkFMOF/++
cFj0G0LOL2H0ZfX1Xp020YkEIwPUXONf+X31gnh/l/1sgzlTTuXupXVTnaFmv/nfmt2aayEm/dID
66o3KezJF67zVXp19jqFzzzqQZOIjcV8J8K4zzGj0eRWiyRYjMAC/WHbz3C9gnvKtH2aIK25euWN
QX6/gyomlYYsoTooit6aObFoUQ/OqXwDtdLa2ROwK8/i5Gfie8NDpLtrs7DrQ2DwY0A/8tAucPaZ
rwUj2zO+fYIGqxcPBFqGq6DpbE4UrQ/K3zjU9elP25lnZ7Jag4Gh2yC325WlDzDizGj/yIIy5PGW
suLRtRugCRj28/Ny9fiFWeHUMvokjUIWNrT4Sfbc9ukGKxtg2kgC6zP4P73hYP5Femb5sztsQTgy
/D7dssJwzOSKcVE/xwDEx8AX0tY7S44e/oOH3qYGRP38SlMuFbbbo36VFVrjjEvUwFWuPTO1MrCO
laZudySrw5VDIxtSirzwHrEDUYa8h21BEpWIN70tLboEb+dAFZsVrK+iYfdW5ZK3/5PoxcNE/hYB
df3/ApA7beNfFJb4bOW12CcC6qVgsIr3wCEgD3MPMLKG3p5I3sOEDbYSXCmebYZRu6NCanIsUyLC
U7tK1X4qr6jpWeSV6Dub8vxxvFaVcx0TVP9UOw93q6g84cEXzR75cvHTQulhsmITJ7J89yb5IXcO
dnCHfmdaFYNyYxw/FqeXCQYqNbvHMJcRtpRGFsucYQxHs93EwpakGvOTtCBo7AaYmSWcRHldPWRu
jwCKyorcvYBHnWPl9kCYp96Bo0OEy36TrkUhGSi2LKuOjvxsy42mySuLO/JesVXfSl9ksvsBKUcI
Hpb6OlcZ5wje2o2kRveSwvklSbTqYhuU5Vi9mePNVnAwl4/dmoAqLscfn3UkhCGH4TmILpB8j2tb
hQ4MM5Wgi1lPcLLftm25TwSnlSXIAuqH6NvpAi7EfBJgEr/3c5rVPR16uya69v8smXE5upd25jMl
/0EP1djrUkf06nAtnMGAU0ItCwwfWWaAApc7nUeCxIsWlvMQ/FljuOnhcOk4QafxN+3qPMJxM2zv
kYmbFcmikVn5UPOmeDhCao2ceJBwlpQkEBAgix1IGdhDzTEmuUNHx6o08xYby4bzCuGmu5WWD9pY
SWadlh2G8tR6o7MxRr40IQ2wzPtDiSP1I3RlH2YPCBSXOzg6bTT6ve5nS9lP8/Tc/uCzacZQU61W
oQl+VFa2PTi74rbq0Mah3IkuJts7zJXNQ0qRSkI0g4RYcyxs/O+YQRLY233dvCtspApv8gxKz8pm
ZGZRmb4OwIrGZhoDoROzNX458imxD/p5zGM23SCgMtOHowUfKRemrLxHB49euLg6iitZ4ZOlUC1y
AdIrEQ+IwfdpKo8NV9Y3JuY8FXfPqfCUd93Ql6aQNrf/sJWIgVLhhXeo85jA1/bErUP0HKcUX1Yh
YiqTgmU6Uz3DzifG1LhgBdFJeIsuGhmjik0LcdXT++r0yIrj5zSS/+pNwEFwvLfiLQRFfSLba5hv
apirkQE+Nnx3UwJkfQNmTaMyO+fjYalKywhdRKijm7rf4D7IkJK+qHdVvopDro9N6rA1VLS4hK2g
jJ55guXFB+Up8H9GLFXnrZqjZBEuWoWz+1miszzZfyKU5NjelGbs+/Wc0B8NJ2+LkgRGlJEDPp3y
CLxUfBEoydwn3rkUqruUe/Uo4gBuDP3jYcBBHJU41nEOKCrr8xxCrOIn8E2HMrgUCFxRZyPFdd+u
+hpz5aDxCEt77slzALG9uXpVGhN/SU3to95RdeM+7P+dNK/g4kNaIkQ5KnhRgVydqh3ZTGgfZbcX
cGP8Lt4UvJ8Bmfs2JgWsLaCcSfge0QQBMTDQFhv9Orl+lPb45XvILYrxpv7KpVhdo1t8TMBl6xF/
2zh+g2X25F9N29pMILRcmTdPIeEyaaRPjiPg80DsanJYr4w7rFJ8wi15Wv1fNI1aEuK/1pXkoYdm
Mwv8VA8jWSp/fps5nFaQbh8Rj6sUX5AbsPr7vr87p22iDYH77sk+Lgwk0PuRwMbt9BagO1o6rAoB
qpauMS2DEshjgUZoBNwG9jbApiKDU59LMaRSZA8s1mx0oIFL+9f8PCLUzjmt7l2NgJpAMujc/8hK
x8lRLystHeX0cwuU3LTAnOQZvl8v9A3oeMVCkee5Gu2KnChFLRB5Y+nZwvoLB+fb5CbgNkG+yauQ
Ud+F16vh3q4tKG27Ves+FkhFDT+X3RnKbGYiO4w6dMrmYy0ouL+e+lOALtCmOedfwAN1s++CD30C
LD/l440tUotDSjwMnsphe2pcPsUJi4NPDR9RoR2lyvOYecE1txqp4561+yW5CTrfo/5ymSge6HHi
HcLAwyWK5kOozeDSStW4DFflxpoB/gdfaZxkCGiRmITKyycTcPDySZzxMq8u5V/73oA6VfO54Vzd
zqxE7QBNO7ZtT1LbLqawX03VCPt0P+z5gJEX3mdNAe/7SxUh6XnGw/LbLiXJcxh6jgyrOBfuWK2V
EU56BCRMYY+CFzWo//YFtStOzzpqXPfj+YgOUE17H6z8qQtFou25ZXIGBXerWMWJuD6ZZwsZ8dhb
F8zofjlQ9fzH14zyXqy4LhV5StNq49iDmKm4lprvTmrhjEqqzzrAXGS7MsqkZqpbk9jM4cSy1xNI
8QanDcVmHf/BbjaYN0lbIVNv1jXjOyLyyGBF9YVoZoRXEdAedex3ecmDiz+4nkhX4YWO6n0fXZdc
8fp2lNyezECIpin6b+3A50whPsPgCuSkZ90oPwDz+1HYNRW7WxK1vRaaU/Vs1JGh8tC5ZYf9EEa2
WoT8xR+QHU44/Zc38r8vidS2+r4/giAyMnfVp2VfpdcHXT/SzZ6rR0/rYPpUe2VWWdp6y5LCzQPs
SlTjgeKmM3SPX03r0LuL3+D0tntIqFlprYOxDFF7XpZrX9OSajfu+lJFi2NHsNYezQOP54VHuzYc
9KZMcj3pF/xIXUONOxs6PXDi1jyekMghBD/6esATz1NaTQyOmFtdxrJxlGNjYf08oyeK++BTCzHC
6s7FIdetJ4WlZk/S1/puU5mF2JvvGqhBuIdH0bIyvpgR1K+FbZa07bQBHMvLwAs/zh6fDEFZLvSd
2kUwAIGigelBKXx08+FEPxSw1HcZsGnTLDU2L7zYrDJ6AY0TjEbsvI3e7MobOkTCVkJYgQVoJbGs
elZobuj+k5hwi6zwrYXBy8ysYgx3/t7Gwyo37Bl8WAsuERAY6pQNh45I+LL1qAbKmtr9tx7qCmLG
9HO3EZ8xD0hcHpFN72DHDufVjpic8QcrvP6dmpSEcGq9cnPw4IqKbJ2aT35CupP/fmSGTxIqH6kv
q4MNgEUBHv9TXShLyRJwzLNePVJ9VpFHu+nITnV5iOykIhoV/KIID/HkjP9N3nb1JyMfL0wxYWKr
rZUYjgNI+PhFFlvlwPzJUhhwyw25mbuJaAIvajiTp8xK7lPqkR7QYQRojxMMky6bJI5RZoXOgn1H
eZecBTj6zZv4WpNPP3NvArKIdt2pjtKwGudhxkgjE1NCjsQk+fWMhQTn1GW56BECwO+VPbP1+hqs
1oEfUILY8QW0g9jNKh9cBgyTODSunFkRPgrPB7a/Mcowq2KYyTxp2HFbQRfuZsAWyNSWafYLb3YP
krP0QF2mURb8E+kKxEziC0Nlyqra8j6OSzv7C5SL+yAScD1PDxLSBOa+MWPdexJf9SxPWtvGgeAG
L3IuiZeNnDtJ7pad0vKXVb4KsbgTzz7S40GD4LCHRL0ZzwUYrBkXWd33I4VDQbhkzarcP3cb9zWb
1d8duhEfpU/2baVKmcs6CGsIs/ehvnf2CR1ACV7+qlIy168sCYYx2bgFQbqxE6aAa0Fa317wVCbi
BTXNtvfLV00dwlWCRkERVAspoUZUl4BOFCDiQP0C3n5Fpz4jxF28CeDIeP9FlXbNbz9copGgl/ug
8HOc5t1yzjgMugqfT8D4ru+jDrF8lOvZs1jrqXqyEl2cfOxatNPHtZ/BXwusZhr+OSNwGfRzIFRp
+Mf2MYKDTTGf4N9kAMflUgaZdwy6r/5ha2wLCCxRJJwfxatuJpAY5/3BxnEXnkdssnNzFg/nolNS
kXRbUYH9eFfAIWUY/Yuyg+JAeibY2NwH+EHsGx0DWmCsglGRDKGo24JECE+LdfPFjGDSmc7CPRg7
bX/g3XM8Cgnu8lM72TXmnYggBsEfDlxyL7lxmSdJtGKuTETYsjpQQCGxvBp2nWZTkI91hARF4gTY
OZ19T/B1A7jQrp9yGGlVY+INVB33gOBAY76wii5OkcIbTIzJMVG9+eyAXLqeti20LIlsK9G1+lHb
TcVZTP7sD0fMqhztLUcZyj0G1IIGsYBjSZd+Ocpuc8wqJOZ9rHK+iPKrLlzRk/V/RQdUOsUW3IIp
wwle5+1FMLZWgE35H/9TNcFbJonK9Sw0gwlUrp6kpIbBkQiEk+sO1rOSdofusN+fP5mBNY3y9rch
n/Jycj3Aidfhjd+daS5Ka3HyvQ7qn7IRGAsoM1+NflNLx/FPdeOYOIJ3V5TrkI7GpsQhtIMEHZt+
rwIJ+owwLP2ylYl+m0tQr7f1xHmlTgztNyYY601lKoH21f0/Pp0X8/IdfFoEtbIldF42WZdqmFDr
FJqb3cyVQJ3J47//QWk7Ei/tXn2eSK3GwAFrzZC4HmKPhGnrK+UvQ37GtkcD+zhlKBfqH1+UOXzN
TsOylu1WQHCn/ydQ1mjTGOYEmdKQcj2qt+JUz37QDcpPNpXi63onrVY1cr6ntqSPlfTMpAooi+O4
Y1eveOYZjxGaR/5u992Nw7r36NNnGbpVGVMWv0nrqbJiem0M6tjR0N1s6nEtp6hAVLpvlzSAyDh9
L61kNuB9UIw7MEryyN4jmYpy6LaNm4wXT+CMz6wQzv+sMvpV1lN7u4m8t3e4brXZEq6w9qaz/dnP
D0iC0Ku8dmD9TlC/igAB8R8ocLoLwwBiZuEb/s+ffr9kSF4ngy8AUqQrGVfwsVgKUPcDj33Bd2b1
fZeWXtkwUN5BoQR3vJjNjI/Sc/c4sBal0iA7v016zFG04c9nQp71jYu4q8bLGQ20cojSIwncJZBC
jWbJs2JhW6bFc6iTbCG3n9VmCDGstJlbYQtEetjlGvmrKAqBlRqeWyGemvSEV+CSDKCVGoT1u1uL
QF0ylNWrAuaoK03ZZjGHbby/h5K8nin+Ue8mjt5hGHLF3SG/txlIxrBrAe8nMxwehlxWBntwJw6X
fgAaVSV3wEeaTYhQprGvlll4ZOOGxkIQ4qnTsGljr5C1vi0FzFDxCzU8fQVYS/9Z1GenI5XTndtg
Zxv7ziYkVoggVC8Su+ID18x7cZnxY8PL7qbMZ3akVMAfAZqXUhbhWWeiB8Qaw/xyVnDTt1UxSYoY
1o8kv1cHLA0NHqstkarMAKuJDppYNiAs3gnELfVu+LJYgQKR4UIXR1mtAs7lWBxGsbvwall5nxB/
3JMAErbk0MXZSuw+zSb6qCPbZUMflYZ9wYtFVWLBhgty2W5yoKKYWcaLPrRrRC/17NvM9tlPUlFh
obMXwcZSx8Kg9YbC2FVqaUyZwiAaOp8yVpcGNQFX6f5FxwtTL7Nq8ruprk8fAKXvn9KMl+u9y32q
LHsuMbo6O+zWnDQPpOD6IcjkljpKQ5G82EPqmjQpuEE0O6/R26JGoR9xNZhGTKaiBbKciafvJNVv
flUI/wUp8Zmotnkik8s4SePbRd4EexQgAaUlRj91DZTuHl+VyN9AZ9bRNQyO1ryLD1ZW/FAMDEHS
n3PhUgdJ0EH3XaeCgnZpzACI4m78IwC9YedTx3YYtR7s5z/0BLfdT8ZUr+YXL02Tuv012NxFtsMC
JyfY7oGBcnVNzf+55PC0xS2sEBI8ZwXPGfUtTahrfO8dxqeeB2Xzbxf4m20x8kxkK5ClqZi5hQPv
XH20PkxjpaNhSx7jQOx38t2bkaMMZt2tCgHWKzqni/zACrI6zwPMADefztDZ0437LHFCc/2FpgKd
NfMSjekQxiMvNBGYYNKnzjgvkiT4pE2wDMmPyyE+RMKqkFwyIwH1OyFNbB6HFH27atfqNhfk6qIq
NKQv5i6yDfYUV3cWHBzcPs7dj/4Y3FfBl5by8vh9m9HVDusmzn+yO6gjSt7bQKwvwNRlm0bgbv2L
GjJHXv/0+6U4v/AOMUAq9i1pkteslDg/Xy8gWdLNqZwQ4E1XgLYcB1hO28E8zG7HsMNhf+1z6rBY
Bedpe82mkZC9P+7IKf7IT6LxypzTnZKAiV/ant0CjZj6PI5WlauL2PMxtALNSQNA7KjV7pjsTeip
rD0bZK/Vc0tz0Nn8e+mhvMWwrZJBJOrpV6XJCaEBGu4ZJdB0hZU7U8fnSMx7ovqk83rzaR/4gQSP
N6l6IBTr+fFgbD5jye4QQdJlSL5EwRKnHnjy7McNwiXCAlbgDCysnr47HvqlJl1p/N7L8zISdTYU
4kd0un+4WuvvA0Y+WSWdwp1DGesu39OyQ1YeQuqtgAoZ5TImOq1kAlE/kk8IVUH70PmO33qBJHQh
JlywfpY7I/2i5XzIJpfN/KaC3rhGoLoNCtvPyAwPqvb5oMlRmfra8w28iL+IV1guh6dlGqlypopj
jJoVKt1tzcvST5ybM0aS7XPUYIK6SvMjUnqEyWxaoKkhHmckloH3GzMG+btJmvSPqvZ33+3F1/oF
kdH0zDqXpPJfO7Uwx+/yMA38/1c/BfPOmoZ+AhyhuJG63t7vrXf+4grQEaMWlJqS4M6VZ+oHeNb/
lr5aWVpd5FZedPk567q4C2jpMQa5+7LQqqT0gIRvzJyTMiIi3Ck4key3zrSQrSLvTdR1MmWHaiVC
Q99v7hefzCaCwaYqHZKyHwsQKaP7xMJfPuieSUba7H1wKx7mbNAkRbIjhgSKq+eXly3NR7cU5Mf+
D+VGlIqtnRb0KIU0ft1PuQ/5nqCBqnRk+pTAGdaQAbVO2QXpcYRcxKwoB25SC+ot1hBN+CbhWatO
sLWtL3wfrXo213GpKe7RiSZvyoGnU/cGqOSmxVEKAXqrm+/e3zKtfe/8OVBKWf+VKcRMp1EcQmUQ
GGBMr6HepxLiM7aotpDMRlzSFDYDWIV4KNYl8+K7cICDp99k5rQ6sG8hCd4owZXDBmRkKC1hNtL8
KFhx+FnhGsSp0cduFjr/ysxVlNX6hbEp19XYLyjYv+8rfXLXUF08wXYbBqVBNFUhc+CUDIUt6McT
V/6i5BQO4GM1C7s7yJuubfCzV5+bP07vWy5Hu+qctmWPa29oEpccPnDk8YCtybsF+SKgZWzMX571
kWBsDi6WB378Ov+bsF3xfn7RWXPP7pDaclb4a7uBH/1WcKqiPNcyiCZ/nF0u0xtOohT7/J15CqWp
BcgvoaeSN1RwPqElDcnnLDGVDI4NtBUxySZ6jKZr8xF/fAv5VlOZI1MCQRhKkXskuMQsYhtr3DrK
JC4PC9pytsqhQ3uhfrKOC6MP5MWjVFxpw2qIxrAGwq4ddyAaX+cjdK4KUqAyJfN48O4ASQkuhpT7
/huEdBj5UYx3tymgORGT2uhzFAU+YDkh88wNIsqa1IPiaacE9MxIVpKLIxpEiYF+BPBW7o6xl2Tt
Jvutszij4DfgXZZkpbuB7sX5khpehWqqDky5Im1gLh+zGsvHiTeJ57303hNs7N7GcNZ32un7wbLZ
YBDofYrkdwVHn0eY2JYqURNMh1aNyw+ZYwtpulVm1p0ZFMoZYDpzY718G1qbpuEeNi4+Hifqy1GV
F/ZRogcouBKUbQPp36dgghpBTfghqEJY0E5bhpzS8QBH9yykyUwvl8Mrzc4ynfq0yajg523EPhz8
H4KyKNKGD9qLvBsBOsyRmiciWECIJxZoLD6HtPiLU1RuYietVrrO0J5EKCJhxX2FyFJ9IK1jfttW
SG4N3+wore/edoguGcTOsn70/2J//DeqHYJ94wRgLgQpEGuV5xLbAMcmH8TmI0YwkjTA+4meiyqH
LpEZVSCxyhup4XGjNd8WTV6n+SkrWqINkjAUJhR0AbQkjGnu1+xgbJhcQvEvypytCAfVzcqk/VS4
acQs9SQlk++HFtzp/Ho64Sh25NllTnYO3ao+CdqxPl7PAeErC1QqkvQ8W/j5FA6wpTOORld2bZwY
4pWKMYYv+G8udbOOJq6t1WcQqX67/UU0TxyIg2zYrBEOmETF+G7t3ZK56rs4ngpvfWP8LLrfUi+R
VpEUGz+DlODZeyusWLGnbHx2jVNejSgC81DDJ9a9ULrTm0zDeie0omKt4gxrFQPwi9kEhPAYM/KD
bqBVJt1Hfh1XNpoU6mENzMmcGnsdieE0TeJKnfOB20iKCRj2YmM7vAod8mUiauzMvYG39MxjXIVq
fCVCL9r1bOSgmrvxYjzUuiWEYFR8CrwjyNdlT8Y8eknKoMMkploFogzIjvd0aZ3RoG361m9oVMEk
q6RBp1TSPb1VQxaKo6VqquXCF1++WfjV93EJqKHzD4nmGb/MA+Szpak4vDC3XQPGOiQQAguZvCD0
GFterffsLclp350eq5BWFbV/VjruskFrzoATfLnAwHc7j5NussEhLqFR2CGnQC9pF2lIFwCfegTL
qfp41eFMe+LUkdC04K65YGP/T7F7o1b6GGxukvUKTFwpfDKpJSJVJPB57bcnJAPFn8HJhA0uTKh+
8D4O+DU4acVO8wRUx2VCaGF0zLOlNJNTBo/WGl8/se6Hw2TtLAO2U7LjU9nj7FQEsGH03QcYS3Fc
7DmJw+QgoUviEQnfv01u9vCtU3SZ+ZruVu2q2qTY3vTNHWB6yc4Yc5DWD8yRTvNhdQlld1C032di
81s7l2aCRBQkKTbP/SoN/mCy42v/MbIXXpYniRZf8PtNQlpfwoeFjJXaerjKJQqTyUauzt4xY+CJ
z7rLDF84X+hXqHc9/xCOn7Z6E6XKLx55V7uAybfTjHrL+zwWvYrO/Dnr443VmF8IM3Nds+ugERCG
1Xwc3Itoo/VV+IZlvXqXHqSZUyUMqnJWBCmsqtMEl5bR3DZNEdL7QETgXcaim+cPrQsE8RUkAE7C
esHrIT5V0iXcnupRgYmdgiFYsc87KaNiQfwq8FEdkgw8iKeF/P65DYRHWFKPXrXf8bllPiPWmmfs
qb558uGVwHvgNJIuBTpYVRwOycNSGYyxnvHrxUnI8dSoV+TElf4PAWmkutnR1jnwGKrcMGUx2ON7
H1rFzgBiFKeNd1vIveD0YOvx8dK3dL0iFKx+sHLthBmktnn5Q6wAKwfxtRypUDYZEQUaHb4qZolm
qcPLEr8k6D+jutOQQwwetSPra4Xrb4W2nJKFTHonkdub8VAOOYJn1M+RxFcNwX1Jg15aT3p8Su1Q
1/bl3MEBe6nP+MZgtpDQtsiGZj2w0OEgZyyM7vyZi0d/PK6kuYJDos9gHdAvqtDDwbBF4zH+21y/
kRoKZ41AYOD+RUueqEnDXdxT8MdmXxnsbLOHZ8FcscrUvKxvoBlFUS1kdiO7TU759vl88AU6hkgb
9j1pgqEzcHkiH4amIKa6kzqsipAT5Nv61pSPPXN3DZ3HHCJoy3MZoTCdm7kL1a1mc0bA6qXcvd1D
T/ZixHaBgYElsVc8LPUxph5QjIVv7XkLjvRoJq4Qzr1xO0Wdr0KIqqzyabFAH88bqPDVeiXDHnhv
W5Q6vRUO3Q2q7UlkjABOL0cGe36e4/I4ndZE+3CoEV97xR5QBOOFWxRBk0cS1FzOdcbGXFkGkFbY
TyCs8st2UscQcNKLv78go5KPPonNX0KV7cXLsSIAgKo4QOC4+axTH1cRy0a+l1opgBfJJgp/dZCu
ZMG7jbu3DnM9MDOYgthbPWrhq1a4rasgkMKfAr1MXz1bJcMuJ9zaXQlWhfiLwmCjBBanrK/Wvg0K
FI9kXR9RjDudXWHAns+9WLBOz+O7NX+GfOIj8AYYkHy0Lwl4pTn8n3bFH9J/QwLEX2kZzIyyxoee
dEJxRkSMXiIlRP2Tjfn6yQCsftxG8XuqzedBYwqlX/rkG9f8hL46NZd2Out2kQ51fm8xqJnHjV8P
lBh8hF6CaX+bsohvgP3Xw5EQjGcK/IefC27Jnq3xOoET73dYdG00VZeqSrnB/bKi2R/TnVtzUV4s
go+MbrMoHM2MH9V6pTUzuxp4jLurg5au6tC6UvezKbPfpOKp2fVW5pAJQozvxBuwSEFJUHLvKk7D
2Z8cN+7rPaK7AZC3oxmGdjDj7fRERblP2iYuMIyDniuGIrs/VmC+mmQy7sx7sQOkFgIuGAZDEDTI
4HGYq51ZVgnzsJJiVZL1txxDwz5hTcdF3Y9TImz2w7gLPMWwdD0KQuFGztHtYXDnR2pb862ENQq3
o6kpCHN22ek/dv7Dun614eX3WSEuhJyEn6v2Cn/o6ag7WuM7g2UrJnFkEb016ttuiHX8cqrN85fC
jBrzW7YovHV8E50RnqSQBJkgA8WiNWA0FF7IetLmFZFwX0IZT4IjruxPdN4wlkTk5EIV0OAXw1TO
KnBDfsmYXph7EDCOz2bY+d22JaTJzJJCmswwjbw7nMSyfYFV2b28yNoFG2oI9EVy3htUrPP2DlLS
pmIIeFuZ6wJcGvtOhCg0aLUP8jcdP4KtplA2+WBXD10h779H4P/1vFRGEtwuRoJ17Ee0Z5y9d9Qi
pimn5fBs/UmhGQc7aYKFWO+6m6r23/2jfv91uvWXg+rmkZMc4eknpzWDF259mlJV7/62hFD+w3rC
WUh4+AnoH5+tJg7nXQESjzna5G+/WXa1L3i1ya2UcKb/CtKD14Sw2oxqNehlCminRlRH4D6ZJW/B
KLTFUFI7KsQ19kCIAf9qIWIA45uZgj5zMTzxN1ClMNYOqxDYQ8HJxD3JcYsKQ/AQlgYwkeaFT9uf
7Qd8bcfbjGdEMLTSzAsU50mGsVH0UilprQWNrRb8rD4Bmtr468k2zBTbk6axV04gQWWvETIh+Sww
VYFAwjtqgdS8+rwn7QmwfsiMm41EA5UKpf7f2GAZ5Hkp60x+FVQe4r/pNHaVJpzy0DwuBUxDBmIu
OTrRB2rKpynu8b4/l9wL8ZqvcYZtNdUS3EmCwoSnC64p1UJutwdsYz3JjlCBv/cFYlKlRIWXw0p1
/dtotSydrqjrO0sT24GWWVwrKsFq/tzkcu0+Zm10YRK7fPCXVdGZsir7rcZnmnm36YDTnL778/Fg
mUsR9vLLi5w/v3biCd1wYr5SWAUHItDJYVwscncVjKWhQ9MzoSqVndpi0gT6tTtUX7pRtgWSaw+S
tIplkT689nYbVkUwaQqZGh8ZnPObOwPOMy7rAS0B1vyxAsihF63xSLreHLSSoHmSmimqCB+FoxkN
d3QlPXx822NUZ12m6AIHMLn93Cl3S/FG7pN+4F+Hk7C4EXeGGjNe9+rTqM4ye2CjN6hxUrMt/KeF
NgbJb6Ud2Z6JgYNrU539fpcLWosdHpYOZq0ns5+JwqAOt7dEe/zwbT12OwGMvptdDsYXE2TGJvF0
UOWrYLM+UYxsoIV5bJqOqV5CR/942TnPNInXHkyo59Xo+x9POlVQcOwPsuTQbHGKzS0OvwOzjruX
dFJI2V/D2zyYyy9DY4Qw8aKjMTNA5CKaoIPwPCKYQKAYQqwA1rkZyxOgplKHeDKC+5MhQA4hdhy5
/ur79ijdZSTa2yiWg2gVkUSBkc8Ts75XVOMAiaX3r/PYrWhlKQlLH/6pR4COMAj2Sgjb1YFLwAxj
M1tans0pHMhJtdKxP3snwdZ04+3uTtEjhtIWyIc7DUYg0ocit4RQ0nS4fnhD8yTd9YdgGs/jA4ls
trfuPzC0IbnLduX54WXeY5JNtXHAh//Bsa85PKVDGzjjz9/CRGxqs+3Qg9bF8rn+8TZ79PFSVFpV
AstC0ZY3N207Ukg7hkuVeBwet5F8u+DkpSF8QvtKTiEBf/BmjOz/PQ91zK/QB4GiXssR/YwlNOoU
/DgEW2ErntreDZ1M04i07x06AwF3kcj/wJSZ0EZplvbFPye+5kEiVhixtKV8kf91ZrVTJreaXt8b
I+ToHqQlVxETsnF57viT9TptBeO6YuKFXQ7s31tTCyo4w8o7vF2RA4S8OQ3KPKfOFs9sQD80tujk
C+vDU3GnVqcXW/TZONgAPM56liWr2D5xWLQk1louseTc/mrXAmgUhkrVC97XWOBW+KYtT63NMG2L
wFksKeYBfW6WO60YCD6jK9ir6vuPP7Rm0n8AtFfdDu2xKq+GNo8AMCEG/bGiWUbemo131iOPiTiD
1r81T1eoqe4NJfjrLQAM4YEKVAH3JVn9UcgVPjQJR4Lbmk8nxYalpRu/Vvr1ocxlbn2pFYyH0sjX
upE8nwolM0awj7YLOIKk3eB5sGxJcPcumtIvvHaGzTwc+gxgVYEe6cs9ebV2DOkfDchZuVIQYdT5
6zmHj7Hh6aRGdEN/NbgucZWZTp55Dx1+M+O1oW3RlktDIFg/FtzyN3aE98xjPlnQTwec1SxAB1oy
CXU4lX4/Qc/iAG/gKn3Bziqt/PFc51iBoASZzSSz4L4RlSqw0He7ZK+X2soX786GpefmrvWuRZy/
BPqIts5DnEizyiTMpyUErCLsg2vA/LMecR6CU3CpT4xDcDVec57jedYej7ZqHVWwrVs8HtKk1weB
vG/eYH6INUviMKOQFmDBzQq5t+PD2bMEQ0Bb/Xne9DAnr/SJib0/Zwe11DDS3AOBfiN8gNuM/Lk3
7j6WX6/Z6sPD2n04dl/d7D78sw0KLYx0jV6SQ5zPsRit9yG/rTRBLNWyrpzykwARdMxVE4tHq3bt
LgzNNCotkgrRfgWppOtDguVLGB8BcGCNhZU+4+uZ8Gcnon6RsD7Ge2BpEdbaW/kFm7AX4D9PSy54
QqbDcYdCOMCAMpgeoW8cFp/rdQhWrij1WejaOS3Oiqyfw3LexHy6A8acCKHOfJR74tlCOcetzh9W
mkw+OnMv8J8MGe81MDGwWWwqzNDQiB86VptODIqbyVLMTzqE3DQYkiVIfM9p2kVjOhV6j2zcP9Dk
8u/rnkTmtHAuewrcscu93UCZbtz4918tL9z7vwpNZMYxCzm2FieN6t82bt6rIzkfhY76VkibHdf3
nFKZemriK0u6ecpR0WfZwv1hBZliVZiMCtMWUfm1oGRmQYn/rpHN+jZj82/iMRBEXDH2It7NomRd
s4LlKlV4hrpathrtMnP5mqxynmA0aio+tBfdmVayS9TA9WZuBU2s1L8aXmxUS5ZT6KgOnKtMiSLC
9i5/1d+YvtfZETi0jSlBJPlQjMa/XON5gN7ED5wkSUW1dvAQHLj/Z95kNm+U8Kv80gkhq+luFe/4
m15aTHje5XPpaRrUkVYo0F4CVxzhugBonAZiANDMSnfV9vpEE2dp3KA3LI2hUKNNVFZFgNUTDSfc
YyOHeL8oFPK3Uz9SVbN/sclE3rSMZNTKj2n4Tw7bF2RtQhVKaj6QTxjKgdBATTbVSmXn6sUpFuV6
pPOyFJl9/zqTyWJqVt1btVG5Cu67dhooogEgohAgjELe3JREHfVoG0MXTR9Zs5pQYg24O6KqsNTd
JrmhaPAWMo6f+YGs+wt5crQ/ZGMKfMeuZmkhxS/DXZWrX/DHnSGzvrfaxlwwZ8FvEBEOd1+aHEWv
Siux+JgOm9HeIOoLL2MxwaJ7oPiqU8DBweBVuLkapBNC7apgqo47kcTY61DeR+wfKaSK8lWjI9Qm
5fv9bayBwiU0ZtXwQ5ls23HngMvBqWsu1Rf37L2D2F9v4nVHK9YUfuLgYhr2QPdy+gJo0mcF/iCd
w0R19T/xhFZK1C2nl485at+YGYPtKBOK9WRZks+wPDxF78/8otedxf8iaNtzrv2WpO2vYeIT+4rm
4LPKzkmYnbzn7bTIGtMrnqZH8/m8e8MYfPVkrVWRGgOnVgFW3GAnyiMCCV7Xiu/mdPAgHi3XmA+L
VWjE8SvjUyEDOT2TdTZhcCEw5Z5Mr5UHuHV3cVK4BtCpsNpRKivG0gYFMbb2oE6uRQy3dYEFHF+Q
QhJMsg/wKtXD8tCjrtDN8Ee7SRR/d0ymtRhX3lkwhpDvOoTkeUZ65mceCwGx/xM7/5MAjPTIkoll
p/NZQLszmNRO/sGHjGlEJ2Bsa76vZBhrVVuIwtksL+tSFijbjx9zcxHlpz1NTRZS9FaFTzk23MDs
MjydkIcm499AuBz/qN2uEHWEiEzS8Q1ixsveFgz9Kno2Ax2AspxdUzcICB5hTmJMUYPsXNr36ZX8
gTwZXbDHKWW2VBAmxWyfm7QKqQMNQDAuobsBXpLmBwuzrqDYj59P6872T5EkORpLJVYLb8sfdFNK
fzl+3W3gknngVGpi2zpjPuhWcdflBkwTpxU+i+crYXtj5dVmdRLV0YQ8EK2NFAuNOAGWGLgipXyP
Yip+D6jn+60lv9fesfFlNuK7A/01AuFQqezaJGSHRGXbwYiJrAqsfkesSKoBy9bW8JKx1G7ehDiI
Q6F82gAatkM0Pf21phgVtqG9Q03bcNcrdoGTGi4BfFrzOmtG9LBSRRbzKioO+7g7DFIgicZVvOEl
3myX7A0QlWJzeuqWxh4dgTl7rQkD9MsV54EFfNEYCk0+fB4Wfb34JlJ2TjmnSoqr/KKAfoFvfYPY
ShSwIpSE9TRYbxIez1MbUQwFUvYy8LH+P7SbQPvWkpOxBYhAq8BFfXfzb9xqlGajFKwbDQ8jgy1d
j419cU8DZEoP6s+Eco3SwAGxBV4WueraS0FjilEwoB4+V+oBLGfTXywwf2vr2rXARFUrodlQ/x0+
3AYsi5GTVfw3cTeUNvI0vj+NHZd2EX1TDn8LYot0MfeNhF9EGF10R8PalydYWh6LjlWmfpxaBbwy
0JTBidmLjNBbgjs7RARArsmdvf47DoJp8T0Mx1Fb7ma68J8tOpydDhOMo+94gKBW65hQ8MSVRfqI
OavFUjDe14fkyQ75XIVEy3OojLYN9zISmSpWv7w3snFVZq7Mj/hXMwZ3xnJx7BNYE1BzujbnSO60
r195sa3pTmTGTPac8HqPqrtLAoviRlgEKgm+gpzAUtNq5hScOuDxFDWePkP9hsOxhtWd8PUVk46B
XOy5F1qCRWhKfuE3RhNBXQtWBlcEwZ+Y1tUIeYCpCdFaO8bi1rKmGlcR3AzR7E2PxLmUBXV25+G/
kLrCfEln2M74I79qepktZr6m/DuYVsf1GYLh5+Wg6F2xj1lS/rt9jjByDLTDozqV4XfI0XeIa6op
X7ABjCrMKAMbqEjyox5cVkBr1PIDkqN+numc0ko6YoeoVVo3eeeaZYeQ9mUwVCfPUQdyp9b+w7P1
TGQdo6CsBOIFe+t7rxlaiFhHhClHbeUkmvcQvRzqr/vqmZ4U5RT/dBu8uxwifAt66EiH/22CQtN5
sAWc/LxSN2Y+dSXvfK5MfV3Tm67PYOQLVpIGgyyo5+bJGbODGvpYZ8HGTclPM4kd4IJauSLs3eJq
m2J4WRT6BXSGnFY0ggrCiH1a7ZuFWn76IOTpaA+rjIvHeLReGP7VWaFFDNHMM0+2NBOU9PUBdmly
oU/qxTU17wDrqokrw5+0e512MNVIoZlbKdWQhUZXY2a1Pf76SLhFDWHaEmTWJ8pStrpExkAuWrPc
QIe8gZkAzBAAh71X7INa1mJAUjJUM6z+FcYKH6rgxnmUHowx9iW7vFU9Z+s0PqSfvMPww9fBUMI3
iema8HrFf7Uo3x/j0aR0yUhMKq9aQ7ngRhveSD4IDKWlDvBUG+VrYzrE+TvCyUgu0rwH5P4Di2v1
6346Dp4rIx82qe0Memr7C8yEgwAA6dyJh+peY2ftWl48N53FbxeBEFn3ZIY4he+J8mhG3hNy4aPx
2tLzenu4s32rH+Mbv2Y7FyVc+tz5eapG+LTXNj68chtguxJs+F8tVPW2QsE4LWcN9g4DP1OMRDPm
vMFPrqlErCcRj6RTdItaL/7GJDQXoeoQn/2pEHtUecWCJwtUnr2G46bqvgm3HxymdcGSdr4aXYay
OsOZ4gP/0ugau5xwWhqdq3imjk+gMz8c6EgkluNKlXuTeVSD5EQF/2P6f/k6PP+Gtv4uGG1yQv4m
qRBHulDW550RB5iImv3fR84wmkU2Ed7UOcJnqSdZ57RzRwn1lHuVT6ufmkQ/Un8uSnqVWJGcgLce
BUdOb6yUHK5qPV7NdRDb0SWyU2fAla4KwXat95WVRc4k33/y/gNXrD/fW0IUGnRbiX0e+9p1tNaJ
1/STbfQn4wlW+TPhDIDMVO2+b48OE1ckdkpnBVMktrWK2TQPbI2k1ZTTYYa7/0Pc0gJTsbQ+Ug4J
+jC9thjWQtX1eQ850kcKH2TiFr//xn7z7aBS2doP2eCJWNxyg93Om7Si+no9MEj8D86nqLPmSfvo
JEdHKtd+Hxg2RYDqxqJ0UoZowrW8kfNaEerp1PIy7GTgNxmaYLs4MnMiTgdI9c7EaixCt+PkA5IV
kZXX/2ekbFmP4pLihN/PFSfAOJxlGWjfSiSihCmQ3zYcM4mEzGWIZzh3rhVD/+SPq6D4x3XgsYp/
m9gom/DG5tIgo81A2fnfgqMBu2zrcc+zeW2LjLgeMzVhmVI29YSdFoZdmH6p51B6d5HH21zugJXQ
/z8yWY2EvEmVlBlq3DJkkyNn3UDneqTkcpNksOgK1NCvSqRhrGeRryeSiVJ2fRnBQvj1qTGHVbhM
IBcht6vsxhWpsTPr0pbxO0liLw/ofmGiZHbRANcv3SEcy9Pd/4qxE/bN4LkYcroWLum3ziGKinhP
FrZtFYQNDhEURzC034tJH8XKk7HNzI7dN0wjsPvIJp5BaMtiuYbW2eS3BhicQtR4CJJ0ly9OgY4O
IwbM/RNnDQvTL8j4gh3DBpJ2FD8RlVGwr7hHDJKWVbZ9VMckqszd7mgAv2CyqoQYNYfLx9sOuAS1
l9H8p/zWQpKzyTIusvv4zp2LV1iWxg0/XaGpjMzrzghhD6fCsLEpljNjpDkY8l+8f1CM21LShK/x
3b2d3SQKEa4mwrAfbwq71XdsC1mLDJVB0FQmnGfwnFbWaKqcVpbe3m/1VAcgVAKxpt5ZPKGMtOme
OTEvSdTlNYr765SZVxiKKA9zUPMFVVYwu2RHj9CIDhiZyrqyokBKY+YydezTZuQlwerdB64ct3Ay
+y9dfv6SVein3ErgWPH/fJPMDbWauuCtk5QxU7d4CSngNDDlw8LnUwR+ZdS4dE+aglsJVOiHUoqF
67zzQmoJo0+xiIAgGdajOkzpT9bwUmOO+8dvZ6OPQPdCO5aH02PnG9NsSXzc/YVRQnWhdViYck1s
zsVA9cveFiVvgEqzQewnKE7ggBVilEmV1NqLkB12FyOFThXr6i4lJjnMja8b7PFOWMOLczV+dz4T
wc8UX9/VUyOjW+W8xCLNPo+8MkzOO3XMCe9msJoPvTKBS6WaTCEZE2R3mjtHOjwMUUuO8x/fbS//
/I0Rq38bz6HuROrGasbTypJsz7n/wvxyS2I8ZlSOwtikHJ5a23MBFcWe7i+j5PsIlY75mbBqlwuW
9d2ChXecPShq1z23Rt9wchmdflK3eYAlWHKyIofSslRM7tvM87EcK0dUeqhuPjPZoaazLNtAb/oN
CWN3kcioVFjZZJAreC4oJmbJh/KOwaTvO/caXJ0s5yKyiVmhwhCUVYsLz9ZPegEvg/Te4mWIBpq5
aPmT84UtM19p1AW06upl34PeVJZn/yAiepR2YEQ2/4yoUi6I93oD/68sZaj5Jy/P4joQYI/xvN2X
leCo0zRztzz4GuOKAP1AgHjqqJL+t6wgO8qbR129tl9072oNQPRwps1A6hchqGl9Om0AxKZQmJqh
uOt0KUN3JHKotNW7pdTr4TGWd7bh4BKNeR7qdDXwkwaNBqc/onM2WOeXQicdNOIR+6gmZNO3SJKA
datuqH7EUQ6+4kIwM2l0fsnDVqqZEpQzPDmWVo4Az2bcUma8fhNco6a9qP8mnQ1W1tUbpfBkaQNE
9nDf+tCyHSupp4li80il8LX5aucmCQ65k8t52Ynn8SuhSylQ3C1M5/n1lZJBVOCWlLuaSySLiUgh
xTgdD7KxmT90Uo5Fb9TFwugJWbvmxlu+R1aXBP3eb+S8Lc6EFQFKsRLtRIjZh/T1HduZODZnBFQr
NY3ABegDPYGL0sHLuMeyDW7nvL/qgse+dpv73cC18sf4dzO29H5zob5uud0AAAwyJ7Gr49VDmlhA
btni47/03cDELPTD+ftQP+mM6OjAUcHrtV0Y8Rwq3MzNWYgEay37EeyRyZn/6geUlbCJrOJl4RRO
PpVoRDRBLScbZXBL3MusLRCzKVH9loyQ00YHYnZTW4PrPIh3G5wW3yVAYUTEM8BM76i2t8A4Yvna
OC7HK+AL7EngYL36biN5cq/dLWgrlSsX7jAJqFYgzVkwzgK/49wISBLMPoMRrD0OWlIaWwg06Ga0
v8iRSOnMa3j2G/bBW1mSYkm5lhJ3Rz8EZxTE/GwwSwFgzyr5112rHuV6KfZqWy9+ox0TwQMv8kQk
Vutlm5l2SFs4XfSNKT7zeyuJbr2+Wi9WovM05lXjXn6SWXf621PYoGjgA9ItHCF/PSdIiM0mETHc
x22W+sQj1cWlMnBk1ce0KXMH7+FRdd5LnmP8znVlYXZjOKF/gyY4PspFaulvDk8b8A+k0tjLaBKR
kUvCvoFrADRHwe/h0kg41OFrVqWcC0h1ZGUL4meuw0SLQb3WeTGOqI442iKf+d07HfvIeI9n/Pp9
8XF8IxXP07TXjqUMBVv3VKpRrwiGr3NXC5rciwb1iXg45WkTGRXzwfeOofNP7QNs9Dm18WHI5uyi
C41kXuOwoXtjqUr3c7jS8D64JgoXONXIUbQ2XiMbCji3pE/ZxAplWv8an1c9TJmijbeer9/R37AA
KtH7VjKFHERnxKDbt8oX8V+3hExFwWs0bdkOS8ZPd3Wnus3guSqdexaYn2ukALIbLVH7gsrnkZXL
KcxyMTf5TE+oVcXNIV/BKE5UwH7Lba64sW9mcYN6a9nwyv2ZKtgn42fU60HzT/v8ns+zNAyWYGKn
suVjnq1dFOIUz8qwjhHbaFZuQbp6B8NZ0948NyjBvGjSA3BpBMDJtvmI0Nqwfd9iNN/ZarMOsm1J
ZqV2wg/jysr29bOpv6Tg1xuRTOoJly+umz6FMlFX9jgY3WBaW50MOM1oCBIyRTYU/n29xL/JfIph
H3uouBtHxsOwRIcDDMdXEt8WAW5QwoZRTM9wqIzwbIqMOs3EMS63iL8zke/aIdhl+joCVP3lK7aH
BfFpx3ekN5K+8GC8CwsPI0Vts1abLY5vNcVdEwZH+bDceBSuD8wh/BcmSU/ePrNFTDTfimUU+XMR
NPX/qMMLxbFQbq1Iq4Eo1wz4+0H+Oo6AiW8m2xqcoewi8gnQ61Q3y9HbUfhpQbzdr9PfoNi4BXIO
78bHOQqn057k4heGulbyuZVqpxN6GetdZezlhQzqQgPgIu17o7lvq80u0fl7qmJPCDKTqTp2x7qX
wnvUxBXxsc/wdYwuZZc7pkm27h0NKT2yd23d07iHQs7wLxc2vd4WW9r1p/YF8QIfJQ62KzoF2Jqj
8XtiCYzR3oFPl192oH72hLDFIHkocsaluMDHemTrvW5+ttMBTI/TjsyTkepgcJv68gUSuS8kwPsN
gWJANIKKatw+L5kYaiXkpqQi/qfsuRlCabwkRIMYmOOPIhGyguZn8ifoc94MxLqGH/ktvuzOqRmD
IZtiGCoc/e1JjOlekzOmlEiliYohPyQdR5KzeDiUIS/77Ffs7UFWdWsGPWGpoHnj5hi5vuEHJj8C
q8BeHTZfeVJw/yTtDYldcfA6B/1vWop00WkszL6daAFXrlRW61yxHR+q/an+FEt2cJGIbHJWPnPY
3LNdJnUMh5SAM+sqBKKO8bBtDO+PA33kF2czTtfFFLg+N0KMIdgvFNwH4GVvLjm5CMglm92MHoQH
LP42DHSmDD5FsRT1YVRNnofV8ksxycRKvVcUlgfgNTAUdnYscRwQnW28lpIFs0UsYxh+NHaild8K
Hpb/D2Cf31jOLlVtfPDZrD60CKtucsGPsdzR2lLK/s32rxsi7lSC8FjCfYLOW0gG6FnE7HKjNhGR
BdWAlqOtVfnZ2Sk6hACgNKo9ElwucFjeRz9BEB+WD/rBNUUAG3r5/0mYRYmmNzlS0rW/tcV7+tCw
8fCIuW3vhKxK7O9QthDzX+5QZqb87nfSRN+D7AO5+vIZrP7ypP0l5oCDTqYZ6aUYBfQlGBzjNlBw
L3EecohgZmWBAUdYDaW/IaGOGgrHZcAlJiGC1uBt33vxHpIH5h7GeL5BBMFirm6wwRK/d8QrDt8q
/dHx255FydLU8dqu9/ge6NC8NhaBAeK7+w7/3gypdI29utihZQXMNdUyxw5gIbMUS7izFihT8Hbu
OdDREzmF9fF5pAi+IjRtRKRBQJGlt3XODJLPtxFhtuJw25k5yUQGIC1hrKZZQtVhX7N4IVA46uLy
7Vd4ZeMCwtGcdVHSULWyafGQJVNMPxOFX9WNrobvoGmpl0U+xWEMVOv3djA164i9cvnNaoXMfREg
HtEqVI0VmWO9GlPBLolFUCKcSGsno7HnVd9oCPuckym/u09AobU58h3E6VU5y7QbuzqGn80wDRzL
q0b/v4W0QOK6pDJD+0JTbN3mEg1O7496EWgcZlsrw29Bf4A86qz+11G7DhMK/i508NE7Sbnp18/2
oFs4pZkbeNibR/JcI3kTM58q5x9lnOdLK2QSUe4PiXQiFCuEngAJ4B8oGjqIG2kopSliQI44B2GW
YYeN/YNKo9OrVNPu3zx1cRujoC2AFHyfpKQIIJ5eSpSP53a1ZiVEN8viBQu9oYRYBnB9A+O24kRN
Zifsr+UI/vQQM0PQhIM1vN5rLuRTSPWCd4OoOTsRWmZxLG7NHEDAdnQI2kc/6ZcQFEV5q+joST/A
eusr6yvNfXQtylBnpKNTcx53S8JnSDpiFRWOGElAFreujGRA/rIMiAoZPjiZfGUvvFe3oVBgU7nQ
bw10MoDbVFAjBoWdfb0PzWhqQRqjc9EniMriBYv2lvLJfS1VXcJ0KPIpFt4FMbe5AciU2+uCDquW
B4lKeUMfmXZ6tHNTHhSgFLYCFuDatdbxfft1uW4hZMg7uMyhr5dmIzD5qa67MN9eQLomx2Zbs8fR
UIEmYZHI5NELL9kcyMaT9tjvtQsANQSiW4ma1az123WMktPzivRPp98zkAu8xWUiTx0PTdHqKEZT
OSlvU4VQl1dUZXK0lqwMwdNcifXLkqLFmPPLvnUvlL2Zdc/g5EczXW0UmQyaA9oT86CxtmWkAzwY
8FlqEukbepN581dVbwnuio5xFzx6cGRrtT24mNeXDkg/3rhUr6MnLtHV0jlyIb7bGXvxpg7hSQbM
b15i1bf/0h0a9Vn/DNLcBL3mMVhAV7l+e7mmPHoCVG+Y/ZNUoi1cwR4AsZKSvca/NXPZla5urGm+
lsS6629zZ4ug758f+bB4kg9OEzVYWOtIozK+VywPICNF8kxJmGQRzeRn91e2r8u+ocBytROZ/3NO
e86he6MZIxvhhQWQW9MrYMvI8HkRpW6F5UeckBVLowYrijtl6EC93mfR0ZdqaKJpl8Zu98+s8i8W
BcF4cpShEvMwGV1LRNN+ApkMyUdmzdaqL7Pverx4D+UIk3vbd+ZFoxf1poDyxrDGJx0B4drBjDCi
xn+dt5Ujej1REMc8WOUxWx0JmcYezQQDSiJ4gHVAc/dD1Qg173j/fEwAwJZ58Axj/jcFRzyamzbS
8yY9VYzaq1ldMnIHeywnFq+XxgsQzuU1seYnu1h2srjUgVO1ZSF5vqkMexTp8d2cWmxgxUET6Uwm
ScIkz7YgoNG/1T32T+Oaa5sjDlyIrYuDBv6fGdaQ3pW19GYKn6G/ds8Pe8AJup2OaL1zMymORLTf
hBrrplremAyArKkDSw79q5+OLoVGNhH87ryzDVTSwQmePI9uztUcUTp5qopgj/xLHbc5to22mMfj
gIDaMF35mpNtDs/3HNr9m08/jeIfpovs16I8Ec6xD7heP/FEvWPiocmE3lp6QG1PAf9L5FtC6VNb
vJioA5bLBKfZcUnBaBCIwuPTvrzmyiM2ew8zfkTdRX/1eMQCxVMm7jZgsAj+bbVbEGj92BktKoHP
ihyFYRHMBFtaYl1eRMeasZVkYbjdfDc1ZILdgc/FGUjGHDptfSu/AuvuRDj1dQCgvIg1Z2VU6j49
Y7pzLWNumjPZynGXKXtO5Og1JcL9LhlrC/IMUh/HTV/zjHXXkUzkRbGhqvgh61SP5ZVULEvbPmBZ
rhK4WGbinIYNZ0+YVIbiFNIKt4FcuAybDblSvlgSKCwvZlBXNaYjoq6BS83yiMyMOG9qrmoEg/7p
oxd9A5S2TsE3XuB4USXTIbliY4Ms3DZv+WAPwh7m8izrEzu/TS2zVWaOrAJmkzVL2ry4shuXOgcs
KDTJ/32PqYuwVLfmtHuqV0jtAXc/T/+LjGsKpWjL+pFeA4GVmVxEvF4xp729oJM9wOvOTAP/bk5T
rt90pnY56sBiuOb+SVLBty3ol7IP24RZZhhVVxqbr5AAT/dBeM62wNwNBWEvgHmyWxJLz2lMW0HK
u73ZC28FLHicIoT1ueo5LItXoTHuYdsJhSyTz2okrhiJ2Jab3WETtosyCRi+4QhYsLHNKu7sQkFf
2IvIHngA4IwMK5kgfYh2v73RdxCrnYFckSxNuvtLOxo7S5Nq+tyIhJpMhBer1kx6nZ4Uw5L+H2sO
zbbSRUBRFGhnteFVeRQ4JhIE8WK4/br3dQDaH3zvd7w4QxSpciM1dVxeF2CETVC7hIqWQ9JlZeaO
F9mfwaKUyXU/BnlUG/7UqKY9T85FX7bAh++rQkKutyTvneTCB75QUbvC+qM9Wh7wh9cXebk0qunu
1jOhk2yCS9uJaJ2EIvOOPAtBvUt2dNgzOZt27yPkAhKqyYbn1yztMts6PhsYFu+CsK9WJUAMt6ZJ
YqYqs/so2Gr0nfCizpoKznMOcTo8pbjARvKLhpwOFHOMj2Vq+ZggOB+AWhVA2IeOswT8Onl2GOdL
3fITRTgYEw+lgncJSJR5v/zRFcOhkZcGa5ViIt2giAS1OvoGF+gijiC1PwWdDyGEjUttAOog0bLH
ioSwcXi9CpIIUnrV5C345C9qSeDPLs94lw+t+2r3OspJS4OWo3HCbTWj15cVguUPPtiuKCtMjUeO
ZaKgYaXDaHPkdOiXUCbVJRMM6eLvfRo9ww3KmgSZY+r+40lqvidV45V1h7g5OMOzUE9nWdp193MA
tQO2X4pEc0Npx7gvXICUi/yDOvZpWszlgsbyuRZUkUjBx9GGHaE7IZBvxUdrxd6eJeQ9Fa9v3mH8
vL0nxnv0p0/0z08BS22AqCkdieofkS09AGJG6kJPTO26aJFuMHcp/33WexMiopb/2rp/X4VHGyAX
KjGtt+hTgYcJMGbkL5GBHzWa06geBfuLX3BAG4t9DGk/ekDPqKWc4VoR1oKeF+xvdbcUgSpd5suv
6HluuiN20ge9SCOLNrbvfOcTTeJWPq4qd/rD4lJnRSrQrREoo8YIcfSLFmfh0/1QMzMeuD9cVG/K
o4rDrOdxcKemqpsCyYVdoDYaW5WZS8tmkaNB4I8Uh0pkjUtp2vDwhA3nzO3iYY8rEsCDoZxAXcjQ
IIpUGTLDVo6Qy60XiEiSQWChiftF2u6G2Dx9tTRkIAHXrDehEon+PQDbWQ1X55fl9f93a1WRPC41
FLFkHdbRhHajL3egqDlWLBRZjdV2epL2OgraFIDFri+dTWXeC0BtRa26NXTSU8iNghtjsxFNab2P
Jy8elmz+6+tps4JzoHYWDJYoxqpSBgYs/kvoUrQnpVCkl5U271jmIJA0FpCkZs6FTctfumGX0KBK
nmO34Kvj+V8vt4v5PioVDkPT0Wz0b2a89qFk3ufHYQmlUKoSawU3qQmJd8LwCTO4ArccvLG1tDjr
PVWZKSJdzrXlsLWN4QqZuoM90Z2LJw5pU17DCxoqsffihB6FbFRemJgxtDVwk2JdNjoSMt2+WrfR
p1jdne+OavB2b9Px7AbpDcnZl3WzSDHhDcUNLw4VEDVmApHrmLLVPGj4pNHBoAzAvS+4s1JO4/OL
LqAye4meQVFlpRZYgUrwgD8WCkSo/z8zaKuRBhUPfVV//878IMFhC2ydrdpW7TSqXq8deNjdNNk/
wYvAVBMOdmrdSN4q508xr+fd/9HxQFGFWKOoKhFxaBgl3uKWhd0ibrDAKTaatN4EetR+dO0sGGBq
CuI/7l4RBy358cKU3N44AEygDb1/ddrFLt/00HsPjOczILY22n/BjI5XOU0Z4+PQS2Ucu5/z687R
Q1aW6vGTbeCjBJEUfmjEZ/sbvcHnzOY7Sh+aU52WND5+dJpRI5WDGj1gw7dtIFxHxT4oCAvBn136
Xf+ytp+wZhhwmzHqW7A6MPbQbmrgbASLpQMAwSRVWFpp/UWnMF29VMkGL1rey9fekdg03jHGkj4l
fnqoIHKDsYeoqMmqdhLowrGHIVDPADizBoEzln7y1Zkc3Lu8g5zcUZaDyBb4gzfcHOQCl4mWD7Tt
Cyq4hOon7DPAlnW8qN6AhdvVCzNmXVGnKx37N+A9/hROdApTWvVM17ZjDzRox5QttFFnvkr0JP4j
g9wERotJG7CBo2+nVy0I2wPvLw0emdiqZTApT5Kg+JCTXKIl+dssaIzoLAl79jcZ4Yisu6fN61sW
jOb2V+fHvGjd2N7T9ostvcVK8zyoL9my17rJ8NqlWZp1j122xP4uyHiuVGnVQer+VGvXtYTqTQIp
tuStPZg27aMXBrVoz96eOk4zoC6eiyQZlSkfGynjFsUDjs6QlGMEVz3xP/TSzc0CEngyF+8HL8Hz
P1yZUqd0OCDUvEx451btI6llEH2mu+Gxk47PGTbH8hPMdqP9gGSCpuSVJqUnDt49U4DQj7/8vBlo
RiOKgKQW7Tx3hQBqvcIbP0GVUB2sgB5fIAgetOPA9BIvoiq22ocVv+JbQ+OP4shasVoaze0abukN
py51gsLnIfoTz5x4BZ8YHiko1LGm36AeaghToprMw7mPDpbhchGXhWx96iEL4pfDEdBO7uV5hSMV
wigHnjsPJ9ahY0/2Kl21x/C25t5UsJKEFEa3az3RVFUmtmx423gio9UlISbbomamdlU5IxlAE7+Z
yrSnASjSB/omzknQhR+wY8vTBY3r2Fl1hi/pRobggWtC1sMuxW++1puVJx4Q+O0Z1BvBkU16OEnI
4Lw0bJwJThANokV6On0BQkoikZPFpgDeEgze5STiTerRmdyw5XovaTnXJXyqyt++ZuznCIN6dnc1
y4Gr1Iid8O0E+9Ecbpe668dWDSNjVnbNgm8cITS5JlQ2HvhGibzVOtsJ+d/hO9dnqPQ+Q+Y5Me/M
zkeoek/LsoA7Ppor3XH8+9KW57QUS1FBa2iKIgF2huOf/S0ItANVM29IDawbtkL+9B8WPk8Rb+x1
/+QGnzLUoFAEpHZn8HzSWK92G+kVu3drh8D8oZbmUbZwle4BiwO2LUv7bMUkqLNwkF9EZ+G65xiC
NGIH12uSVwL0jWCfZM+A9BkKF/9Kzsysj022o9rOh/4ltvVsQXOwZ6v+JllujyEhd9p6B/ZfkwNk
tIOh25fRi0ogQpY1bft4b45CE2YUOJqRIH/3PJMw+BKJJteyneAtqWm++IJtSbzHQ18loOFfkEA4
lnVPo64F9SQsWro/Hq5bUqUA9anlDTWUsyaqVfxVMDDiPLpCxgtwuVzwxBw+oCOu6isDT0lzNnhu
AEq8uRnB+bdYmpWsU7j9hfIRTzji4wkJWZlA0dSzy708iI7GFeYVzxKnXGiz2Gu7l4dBhjmPYjif
EuOY06ywKReCaq+afcaTozw0d8p/tkAEI28pU8pbqqgDjNjfdebnlvEtm3rOExtIcEfxGbL1u7Ut
h6FSNj7uYF8osx66z5J+8OJa7AduGd25qs2JXk0E2KtEkrz/AbN5UyCEB5AChj7N/zIaupJ29Lyj
JI/hpvWCA9hd3UGwT9q+meqRJvHpQPSZvwJicBhYPt/UeMEAwzaS3ZqwhF/2ykjbPSxx5ebyOgQ/
phpnPfw7KXVMqebaIvXC0v2un7b+LpZ0AYbX3ERlMKN70/9lCABPyapy3bC3VzwNX8SvCXljt87U
0QW8UhpgVaOqt9hRxn00CzLtkGh5JqenbOcJS67SHJa0ixMfPD8MlJStDE/58fo/jETzTVVDEitH
rHPqz4fVN2tXvLZWc+W+pMB2jwLPkjC1fQ4xc1FH03vZvAEJV5x2oRadAG8dpEVdpKzJlru4lg31
KBNCDoBo61vA20uUPvbzc9uBbDDOC6Sh4XWMg5KGxwtsAm4YsNzFgYdiYJy9xSbKI7wM/+O5+qrQ
YA2SnGo+R6BDP23TMMaelKwPiDl1P6L8UAB663GmtdohvURDRZonYFWQlAzlFheFQgkwdfryB7NS
ewZ/jG4FtyncnCW0oCkUIQsBdncm1SIr3ehaSD7/rQ6M1Ptey9KqxV+mFferol3NYi8YeTEfq3oe
cQEDn25N4Qk8/cqw2l/gyUWnsHaahgY8wveRR82NlbHXoMZmmX6aaVpXzzJEsMSanUIKFICXLMsU
NKnqNrzscFpufyg6eZ0L+YZ+37DguS3WhOjiCusTe0v1XU4Su3K/ZvP0dqTd731/J44Rch/wtELw
eg13BA8f9xAoxCmn6uP7F8r7x3m3SdYC7pfuGR4UQ5PBChMEvW4VTjLMxgNRJqjIJJ1MfV6DFwwz
WB5qH9cjr5ThuqUiekLlvC4KiemfLFwNLx/GgcKopIcuZidBpUhK/n85buv9voBIq9YiE4piQziu
jqpNnmVeAizn3NTnjsGI+0KwUmTwcjMPYBkfHqBsLCdE+5dwRihUHRRqGMg9mIgDuzsnYBh09Wxw
kCWiTJCZ3QW4T4xLRasWwv/cP6HakHZFapd0P4EIphoqm5Vh6xPcqgPrt5EGb1XyBY7Jx3+IwRBk
tilgKGYZhwRb2c3OX0XZfyROy+s3SxzxT6LmcWFHLGDQaxv1Yti0YlRcARUpcU9Lv3kFDJ03uFDD
IXXIrrlcakPjSqY0PAGkj7x38Yd9PZh+u5KZiUIP8enkdHwgT+tkqLaKnbgj2YkM5uKYjBLcyJzs
vTRqFxa2zzaFfcOREHlwilp6jR+5gBIrzht2otbxsPJP2GGaveWJSqiyLMm6MaH1ytdrUoaoZ0AX
OmAOOVI51nGX0RePU0NDwlzR1fAnatRPnSFN9hLaUNQnibprfgmqYy9UYWFZ8NX+3m6VKUE9BzOb
8htnKLLAE7HgUEdSQbVjPnXybZN0KmKRkeFgcwXwD+AkHJYmmtMNjrMCtdOJI0bs5yziQ5vLUshk
zeOckdQ/sr2jcG31o2untrqs8SXt3ioDC2uZ0qU/QvhRaYmetE+kYfK0CfG+aH6sB1u47s47lOJp
7gqzzMZSosqXF5wxbw+eYz8vYOqKX7LGnEeYqaWhSRXq2X2QANktOznPe773TJMMMf2EoKv5bCza
GUFbrCCD6Wy0kE6CC4m4rfRIb2BknnOP1baAwrv6XSiAibR1uJaAX+C95QIUgpuU22dY3HcORusz
iLsb79Vk7hP+6nWANiqEegGZep2IGpz+ROCoNC1LpSpBVAhE++v1FBYLPOqsV5a0IDCA/uA9Ta8X
gQDohdSpsd7CV9e/yTv6SlJh+YzQVF7a+KRpdcax3z4NoJaMy6eZGFWGbS0aE+NMtExKx9ngVIm1
o7hrmTy6UWzpf52fu0Uw35dUbAMK2+CYqR/duiOOmNCQvCw4LNjVBWxRR2NyWgRtPpA2th/giYTj
Ss2i+95//kC5BTDIFesOeQ6H/6VNUgVtHeEjefsAHzDm7SzkdpKROd3JXjVWh9YyHcg7SXE6Y2i+
e+70ryF1B5qHd3XsiFjqE0tZw58UYFvkdC/rY4dYO5tc6I6jM2uajstcHMCFn8PuBrqxpNrfGMFH
SI+3VAEGdb39+jlPpzljt0TPQtGqEiDTRFzmZB5KRnEi58JILz7WlWe9l7wdZ+bRNd/FUfLmE9aY
nbMR0zuDyqZTVNUEPhM8zIatvGOvgEzO+z/SpP9Y0xNlICyldvwgFNYPjjfNWjh6i1+vXwiZo3iP
w/ZAPZg3yCYRulFl09lGhvQRAkwGAHm1K6qHcdo2DyA24bp6cD3sQaZ+WxyAIQY19nv25mEPs4p1
BLg7c7hjeEHSFS5tUb8ErTR5OkRYUpOq3kSiYIonj/XV7YtKXF/eHYoXC4ObAdAesgx36uR7ak82
kSD3ZVIA/Nn1DacrsKyHdc4tgnkiOdhGpSmgk7WWMWGMStPXK+qpzIV/zmNTZxHlpLSeklGFiJF7
WlhTRY2V7IfFZOO/aXEYZsW3pc47h73xuvpQYjIvi8yiGsfkOfbkjf6uTCVtNRzWPZZHoxgpw0kI
GOpI60y61X9ygKaCiq7vYK+GFq8agwRw7jzVlMAcL0acE6Rz35FUaSJ2OYd69Yb/ZljU2Y5qDWID
2CH5fPi3asePNvPkVL/By6y5dZ89wmCk6xSuc9CPzH2PPtJ0MQ25z5ymDTmpF9OEabyQrttE328k
+8gEbDNGLxf4I8cnzFF0jQhCukRwOUZAQ9+LPBSgVsaMlxMyErrKbX+5/mRrlKqBbKCEAPFpryZW
A7GtaKeXzOAKJG+Z0sgWlc3WQjJPy8mjIBnS/+qZN/vjHnWwlaJUbVVmd5J5khPzTebh3qBH4clv
Y22B+3kpDRH/m+BK0n3U1NdLQh9X8DXqZujWh9bJiNrVp1n8QorXpx5+zj9SNl1M7KDfz1laXBKi
1HuOprmKijq1QWVyUmwnRZQHNsFeVTwTHi9DBJ0oxy0K/qmVtQ0u9/v/gSbz+jwyCsUR4UZoZDBQ
CLlY8cqJ6+qcCm+SmKU1BlY8aVFWzl9f0Cv9x+Qdb8dTpB0l+26DohGVJskFvMPmiqycgKJbyr/V
yBPJJCku5qN3sXDdhbNn1hBGtoe8j33WIyJFdFox8fWEjbqnAu4SieMXChwK4RfNiEduusn7GXdY
INO0cF5PCfQdNcS9osWVTxhBxEAIVB8AM28uSkmnooctwJh45a1BLTakG8wTmEzNkSL7z94yYGd4
NcMsQzEWaeodOPhWpYhYGRHK2oS/3Pg/V7Jv1JbqONxoWyhPTJCx/EJkSa3vnSjcaX4LYIgm4W13
fvpVtSNF59tcWb2cNWjIB0qscBgMsBC+A6dtO/AHtCnmwEqxmrfakBwP45wr4i0ytJwDrC7QOJV6
ctSWjdvMjNKV4y1DZ6b8GUDbI6T2qgxCzAyx1pq6h9WQhPUerk9u4eIlSpxYmcpRQuv8VZZKQTXi
yj9l5Zwdy88incrEPgDkFJk+3C9GWqGZClQ08zh3oxaMAfMeoSprdz0j7BEGDGaRMKSSD43yNGJa
pLB3q0p2cVJq6wLHjFJAaP8Cbdp2UetrSyXvfOfetNQ/iskWMVC/EdUZEGMJ/M7mV/w1ZvMQdE1h
9eZqSnkkjmTesPi5QCkhBDIm+QvLBq/eKrMb67hM/HmoYB1yAUYhXut/OA8lSiEOCrISmwvFypA9
hIuXD74LRYpUTKhBkVVjO1xb+tG4j5wWgRY746aUViY6KcPYNYxXzl8hKMaDoy2pSbf7w7CrXGEz
xvpXpjyE42eZcGxBZBKEFz1DlhnTvpDG8V4XLMQ2UP3bcMW40oK3WWzN9Uw9NHt3PV/yszAFYw/c
u/IqpFyuUPyZZXvQr4x6Ni/3SKSIjdqEfLS1ZyH8LcGmx+Mg2rfNyJXdod2NxcUTjnKq2DkAlRqI
LSdUf39Eq97au8P0h2/u6sFjkeSLqc/2VBtjMy40AYRSqIHVS6v1GbOoPFFlV/yDgC1KcpAAClhO
rRFpA8paunlg53oQ65fNroRb8nTqzhUst9PiBKg0ljFsQ7iAylUgHwzFgwx6TneQR/YXTgrrr/0z
v0AzvHbjBX+eFDWJ7AVOiz8WujKbk1WgxOR2ovlwby6vyj2DJHO/q6s7yoLRPUnYX4X9zlQLYDxw
q2m7luvSiazbqbcGggtihxL0McH0INbiuk6hlGjv3QFz4ZJ66Ytg6sxzu0328baWXUTKKEH1TEL8
o1fHeA/ktI9FLK7ms2rWVrbmGXdqoIbyEtuxBlHKFiKYe5piPTuGYR5fNpm6dA/VNybba8Sm321X
+0y4FlDWxj3ih1AmTatJ20Dk4c5tyuI4QmM3U9jdhF0GaXJDJ1b5rN6tULvrPEe+SO0+B+SELcI6
L7dkmsVXy5hQYb+q1SSQ7blH4LR+dp9S3MTq/Aa8Uerb/1jsOQECh5TvAfgWs1n7ENMtbAZ2hJ4k
zwWa/6FgfoEQgloMp0WUVrYcx+1VmXliZDSvzS7SdP9TuUB5ffW/sPar0Dzdcg4O7hNkUUiLkIWx
THo37wyBbX0rZK85FE5oQ9twBu0JjZ3Bq8mBXTbaZIuR0x1UD0RXnzBty7G4yRgeiV13B3YUt3rx
Tb7H0l4vKjJFwsy8dbH/PZ+x8qtBUykw+Uy3nWV8bEkVCmOp/82ayyQPNmvoBk6j7741V4PqM9vy
lZTgRKs/FCIgcfcmgEk6rLhJ8AkOBiCn5mPV3OW36esdNIIEwpAjitld5IkahMDenPyUqTN7w+r+
LcaN3NlyIIpOi9whMY4pGPcYNrexEUyqHSFPLpASihPV25gs3/4ZKLAX+YWbcY1DNfXcDh6la0V+
+5/7EK59mHkVlm2lH37q4QhgYIHDPxnnJn6rUhY1Dvi6RuEzwcGFhjgNCqiEVxA6bS4MjeQqQF1e
bBEBSya9nvzmop4En74lqzLVJ02kCH9sGEhXwbLo7chM8s4YFeGvBtyRsb3rwKsIRlUJEy3qfNWS
s50zpGkGbbxLrWtVRufoL44POWdo1o66PcLpYHKZNtwVN3G58q4qhtad7Y3nnCxYOF5QfblmmqUJ
g8h1de7K5LKFNnfvcYAAvXMCNNsGEkklnxFhN1/vG6gZebAbCdksLvUXjal0btRLTkZM9hlvVZ3R
1s5XFWzWp6bVerEx5bLrO6FU3BJYvfOHrPNXGyaRS9VuIIc57uuF27tx8WTPvODwZSJ6wUDEyKA7
uuvQOL8L6DniZboyTzil813rPqclGyJMdjYyrSsX1UxWz0x3FOHTDBUObTLS3z3DWSfzllHU3NXi
UBOnbF3d19k5vMqamC3uqve8bfMPB926f20ttOWPen2QiootS5UR0/qcM+x70sXvBVCeW1quUUsk
41i3RLBhWkNMtB3o7YlWDmK+AYD/l28YjhkVnODCi1paw3x2ntI4eEPy0ltQ69OT1qIscjQPo+b/
0Z+mD36piIxdADLFfVtphWDm9pWibwctHALIu/OqXFGG1Qxi86/20JvAXj7iRZY6sDnWTIwMMkvu
QW49Po6jrUpzRehQOXYOVtO2A3H7AqlduLK0KAzCvvyrhqFul2y9Cla+ZjdU/bEtv5xA3As3vDjp
c1dSY64qOV5rsstZQkZKShZl8JRgG0hkFXUnJ7lsl8hOBzyX8rX+mslw3NPT0pt6eVI99IHDd0Rh
s7TXQXEDvp2wTsXZkp2HXUyM4TXBq6FcFZ68Ae1S61ElN9payziIAyVUFNLTrnyZy16uJuK/YUtp
KZUeudeknte2ijqib89NPL48YgA53wP/fb9w72VJYVXgzPD2mGnkFKf9sNX26hsxnM8sALQLt5gE
cB0hK0v3QTCoT3NEyBQQafF51Cfg5Ho/dLhFsiZLWjPCep0FAqed99AnJZ/TYHjD8o2v2wGFFshr
QDD9rQ96CZRDws8HZBiDmkJLDY+uNdouPt507Fd0AxN/V3lraI1foCS+XAEI629glsaUPt3ZRDEI
Pi4aEdNgmd6s5QACPrxeHMFrv1XfbDBLAyQrTyDjqTUssFxI0HztVMTDGVkM5nqklAm4dw/WxN1y
BdQy34tVec1kza+inVVq+LxeEVV3x6MgnHLLfzFmGeHug5HhE11L25j7Js+9aeJ9p38OpffMmyYJ
+JAC4L+pXRyw5XGzgpve564EBCEJ+TnyZExYhsk50B1hn3YW8rCusN+5n48hwXPm96/+UOJRN/AW
p2JKcS0pxI6BZHEqUEnykd9RWoD2KEzyL47lgtWB66Nm0gMOCx9uKx7TQ9sCrh5ElugG8T2mTuO9
iHisLv50yQhPKC1LKE59cP/99KPJkiylese/GXQ2k+vQhakJFRKcPYtdTTXSb81/dVwybJqqJJia
9K542AGGFNoS9O96s4O0Dbd4gMHXJ5Ru6YkEPSUrcIMeBdDCIP3MXJySbuLAnn/UN9XExhKpenY4
QFgDgyzPkim+IfPY6+EWcwFJnldB8aPADg0Xil8pbx+fr3E57qil4DHtqlyuSgQ96iS0nKDmDJPl
bfP0yL1PgH2vtIHv7oDIOcCOGNrdk7QLaZX3uPcrFNw6c+IlrxZYmjFTyeYwxnI1OI44X/YrunbK
KhK1HFQdsHtvhQPdBRKfsHyEsMRy2qrXqowoou6Rn+TQwP0X7v+h9iq0q0Sj4Th9NKUQObOc2Nrp
K23YJm8kdAZwSnuxx0kjmk70YrBE6mnhbMm9CnJhgLiDPEtgxtbe7r2AJqH66OR0fwgzf4UUSsWB
M/msW454bwTCilRoKmpbd5Tr/cVge9vV+Xm5mYqVx3EXyqtOjd/AWBVdImYbCEUxhTEUeJi8m2Zs
CMZpmSoy0kDS5cSaEGVlKxfsn+gS0YLEMHiDhewhJUJXoUFqZFTXrBoc2gwKV9dK6376luKkx6Ct
9ts56PxL6qq/2dQMbtP0TzUt4qY4OV02/nsXILUiKKDve8JA30SIz8OL+2zKkl9xzrnIP6qUYQqb
Xj918RuTj0M9nXzikLRWMz9BM0l5nCP6IeoKQwYfzvukpTxOF/5SHYSKS3XfdWWLFSJq+H0YFQyO
ORG8CJEb2LmaKX1JZGjA1fzdN6tWZ87SLaXb4Tg9nAsK3N4zvWmc4kUhZpryQXkA/EuxyJjT/Grx
NeXvCTf4tct3by6f8P6Zq8YmLgKDHdbjg1nROBmaIwD4+FcKNIP/hOyZMp9Fs6Aduan7bnyHnMqY
ul6DMJlbfaCcw2jPhe9GMEcNQa7llU658fL9pCtk1jJRU8oYPqjB6DWVoSoOOLcRLP6X5haQtXnn
J+NBJeHLFkV1x6m6O0oe48IdVHbyBFbK9G572/niUJEMTZXhinI7TDCBRJtXzzOPQPy/ck11O8Bg
YDVWScF+91xMAIs5TbNg1Y142s3RmcRbeSr/2yvgwPmmRw6DsoWjvOuOCWd1seoPvzJzmeqh+2D8
eISOngL0togQwlW9caoskA3xaKNttnu567Zp+QaiNUlcC+aD+z1YFCPi+ZxbwrBI6TrbXGBF+hya
ceX3m8yb+mD2jki+ygN5w/vlj2a55v57KEs3aAKV6Im5CbYJ0gjRDPBdN+79lHMgj/Ut3olt43U6
+gjO9R7pSkB6Qb81tQwjjDhqEXtHZ2puvkIeFMDHG9ue/zF058/eW2StAd1Gkrh5fe4z4E7KZAX8
z6GX7SB0CeUNx80F1xhRVjiwOGaReyGdQz9JCYltgYMNPa7WP8g4gX3OlRdVH9sKQDtRbCTWFLZH
jtUh48+XrD1M4mxtxzPBbmy1gqahd31AQWmQYIJ0A63aN32w+YgwwUrDtmV2jMicTP7x779RR7Z+
6HUr9Oan2+seKV4YqxPVK7sxPkhbo7w/YsM438ozmTVPK3lKo8Z2mdOUjgzmfEblWQWDrZ6g9ngz
8FbehbTn5AWUv5iphbFwaYy2jRO9jk+iUvN8c4rQ5ckCv9RW5PIXNqGfAX7BbTy+SavSm5jeNJGD
s0CjijObPtyruqFeYcaxnMsRR064TEuUMOOS4oPV3MXvhHHjxW+wTr60PExdNL6WhMYJRdl3kD3Y
PATQgL/qqVsWutQuYRNZ8qvNgl0VqKXB9LNYJ+83j6otKn4ahPNX/HVgz0nCWHyUcUv46X2ds53H
Ilb8q9FkamZI+A6bvNbmpM8bh4vy4HZGtE5gh1tDZ2kTYEDlZCAaYJ7V//n2zDt6sUphWI7QOtab
Sko3NaGv0li2ay2aYnCqTTpjX2Iuwji+zNh7eQ5hgrT53cw6CIFGX2HdIkV1In9QLSwkwNolzF3o
JTaUEhbs0rrcU+z3jrIku4scVUdc4SCERcuDzNe6YoJHPoTNHLwE/H0o7Lb/7OwSKbDiMkPlhIeV
uSgCaNP6btCJMsl/wIKIBZTpQxS65rV9ql/Ijj/fdFmq2x8gAwVQ8pkP2ivh5K+XD1Bdvyd9DoMT
C838d/U5CcVO1iwbIl4UWNCbJL+V353pEG9fVq1+vEmv87MoybAXKZDOktNP0x8w6ZLTEWTGETlf
ALs0R5JCSUzv1NCLI0GSDa1QVvX0w3prHjmaLPzXFsDf6VtJqq4AS5NpuEpkZ79CNlD9XmcZgfG9
UvtBNRl76Q7trRwlmhdSqxrMsMLNQPpyvqRWQlgIUHke3NGbri5RO7cg6P7ttemVC9hmved74ehg
MPEnALErgFDTfl08eHI+llVPEdDAj2QhhDb+wg/BQnw22qVlYEXmL2c1mhRaz8vQc5cqL2kLhnp4
O1q1t/lWbpCSkEVaQB1WCP+Uld96SphIMMwtFLz7lOI8q1rn8VEresbkTCF0/3fscFbE2L4/HhEL
tt77xfi7etltmRQTvZ2lc35DzhJXbT0cuEVf1rOq2TAzl63YN9f6N3l8a+vfytiP31H9BgBi9RP5
8CXIQA19gCNoV8cxDss8i7zApB+wER4ms3jA67XjiukLFStcWm/xHHxFRDiqlh3XjHkMEvutEJa+
kHd9Dd+klx2huywj36DV6Q0q+V/G2GALkyL3SH/fUQS8Sk4BVCqnoUx73iuttL321LD7oyTR/eqt
7/Yvwdl0Vb3f6YhTzQceERCywZdaHqtBjK8VUSMd+VWe2p+jT5xOz8fJGgbLvOjo6+asOTTBvxaI
FMWCNRtXej6NILwtMBc1Leg7OqB70fIzL+t4XDIP5X/XihFrNxTOFOuI+pBJgnkn//jZdAL30BT7
o/qycjgVHXXJumrOfm7WDXQr2y2GKczbFmThfmk1x9nos6F+T6p9oOK/7URcIvd2JRFsUzsLj2Ld
0Yr5BEnqVcUmUuRzBP/6wA7i+lBG5iuXMakxUV5Iafa0Vku2Exw4mUOjwTBkgOUEzbAan1qj0VkR
fcrnROzfbvCNwogHVDq0aqMOEkYFSFq+iH51xHjHAxsnk5EVkPjvfd9N0frpEeYBvgv2meDqHtDA
ZZ1+MCzbFUWeJkk3zRnz24ZRPvphcmjAZNsqw6CC8jJtT8W+JdOUG2bBXT8XNjYSxxM8asEh5/T1
Azfot4L9qzRR01mUH58XntPpzbFP2F10oYRQsx46VVVGjNUx2C7tcegFu0ATtaZfE0N45Absmcn1
1/eBn6SkCwxqpNCm7h613sGyrObIhKdbiTZHBnpWkGdkiFXH5BLwgzy73JkzTuDuT1d5pknfhAMz
iOZ/a0zZTHMYzSiXuPfUoxE8C66YiN/wLGlBIPvtKoSCd5eRfy7j9CyrwW49td1AC+fPaq3SEKoq
TAHnOdMH9p0cnu2evFkTsCqGn5L0o8bsZ+cfvYVxppCq8n0E6lePelLjOQ2+Qr9eTD+UCTp8Nifb
H+J2vhKwVrp3PNNttejF6ThhsXn80CyCRkazFXiK/yme3nfSZLRmUueWmrNElW02f/C2tYJHz5rj
FGJ5sW9zslMW2R/LUxnv/m4oyFnE/yqy0qIoqKK+QoKsBiGmlVSed56Xo8DEcCKoIBYpO3V3JxiN
e/h8X3JdxRMNnurLlpXhruFped68b2zTbuwb7Z+3ZbgKxN3dLjoaFFUXQmPpqXPp8De0tKP5OIrj
Mm9ocxoCegFd68mQORrdlqODUjkhJDKcE/LEFkGUOWx4KHk2M3AMQgZIv22ccF622M+uKxYOYqXA
ylZVirXOE+ID6EsvYo84P6MLdF4SRxMsEPAR3oTug3/fubzhq57KhkI8viLyCJTghuNbgVhCLx2z
j6X2ziXRvYApgxn1hIPAZCZnGQaoEn+WL0UC3iIhbiaI1RoesRTEIcDD36Yy/liWWfLRLonXsSlr
WKS8E6Tqfvuk4SGYzhgSBBWJmqij41HDOjIGoTYBKlkI2fEG9lffZsRvVyMrE0sx9705wNrRKX08
l9MHRwAHt5WivQtBnHTFpIFFXWRAxhSyamA8H6h5qXyZNE/otH1PCv7EbZIbJjwHqFpW7XWx/mZj
ozTUKBKUkTPyojA1IdAidvyLqlosADymjznA5y8nI7EsjiIXI6PzLCoScaKTFpwkfVlBSUgFXuog
GHNNTjEMjxxoB1rgx+d1hlQPL+i6AIzIrVrJmtp3T2atUl0a/wwnSbGF+z8MoEIvU2nL/itQV1I9
omAW+6ydSZISYGzOhZv/OZ545u0E8HqCQ+ILRmxG5ZhTE1bGJg5sRBvaMU5fDFZWi81WIehzrfuQ
IG1FzE8nVpxIIwqoMkEV8E2QGBjNl3SeuQTc15QZ2rE8/DkNRLsBLor3nPRCbptD0KJUA+o/6N4X
mT/bPP4L8+YOsP46hMVd0/Xsjmp8tFucl8mvvT2P5J8Cqff34Mg5VgA4L8CMSczH7Nq77vvuMdrm
rlpLqYdQTCtec2h73SvcN+vKcG7O4tpdqLTDxQUMt3L4L4cZnfdKbq5ZtxLrIWrv5lkv3a6FSl1S
KVXLIFsnBz61y44gT04uFZhYAJQqNa6ly5c20+QzHjRqGcAUzBDo1fHylrvIIGXix5jzytzn9A1S
dzEz3fUDwIDbxmg2/a4IE1B1/ru8pD7J+C64Bz97pznjyg0ecBiDy2HXt1+x+tYye/yQDdfr4efi
2i1yGZJT3/shIbs7Xuz3g2Ii2iI918knW8YnJlJI3lMwhwIFzmCXlG27HfqpdvhpM8cMm3mtxuXG
23yHFreSYE1XDvPSdYL9MzaJnm3PjIUmP3Qnwrk9xpIFAVJ06KkiS8zuDMgpnP63XAyJDGW85chj
kYfXcedcpOPkesXzw10U67dzL+aR7+BOxYVrV/VTKxv8rLzgffBBF2NRPPlXmv+f52Z10l0cvlXt
xtrxNMW4N5rsFLmEgnMDU/ptaiSjloH3loeUE/12EuLLb2XoIJcoRirREYQ9NPXv/LkztFbyyFWJ
ZZbxehMGo0wOVzgqNDknBppa7hcj9RDZWvxo4V0Ogf0akfmfFcsv1KLdzEMd/wHxXCXfdfIfaGuL
P8z8M9V62TMdWdPbCs6lZh7Wndo5KdzTOWbvDofBy6du5kGKU8uZfy9tKkaO4GH2+YjcO1n/Dyyi
HXgY9gahJu3ooVa2unsrOOiHvx2NhMbsXPOZ1CADc0Ay0QNUMsnRQrtG1dgy9g7nK67GnhsxJacW
Dwq90e3Pi47GTBK0obsYVFA5uTMdV9fkAgx6c6cofKhwWQTN5LSwbFapi2mbA4snGwKxBD1M0Qhq
FiCH04RUN6GeksYLcauyhJDe192zFKdTxlCYgooSidTmebf6ZlwisXU3LKkN8BbRhrHgDHS646H/
LfRxM6FbAj3jUw1x+kjLUw0/tdV1TkA2btX1LELSbW8zdD1GjdNVjtRInHYekoVOVt7IKURnVpJL
gMCUM+BwJxZeWBhlwmPyglM6TO28kYZoYbbhs07YanHqvDLEaNaK9zbtzsMdNfpEOVPctnnSFHDT
7cBVO3X7Mq+LyvZuKSwSKQe2CR1dw9K3fLL2M7L8aYRJ3B2s+Na4e+BHy3nIG78MiKdMvdyx4iyu
KNfrREIyGkNTvWouRblvormnqh55IBN88txm5jTNMcL2ZZ5K4z3Mpx2I6W1jXEyY1AK0TyYhPIuj
wDswK4lEEmpgGwtp5xyToFNzPIDnVLOXZxJEWPmjFI5GOnK+MVTrTHcGKmxK2EFHS+vgcW5h3y6f
V1IVOp7VK0iqD5z8f+ETaWePGH2BsduMe+dsIB8kYj3IZitdQCecpRQmiEjh+lNNCgXYvh7YC87e
WXohqcLGqCrUU3l0+8to8XlSPn+yOnloRlOyX11NKx9EMXvvTGPYKq3sJmbBmGkhk7unOrrhK3dU
aTsG6Zwz4k2M9mx2d0Uplo5FdAZiZl0zqmKFb8v2aPlGITFPaIfxoZrocJ4XH5Yc887/W9vPla3x
/jttym+FJzr1X/VUzY9p5mV/z5VtvBedmvnJijKHn7JHZDBhEGbCqpQF40JvlKwtyPfIuKkE1kGr
EzG6ccCGtzKhJUqVHdoX6t6AAvrff0FO6lBl2Fr8Ef16yx4sfZC4lr4pcWHYQtNLtzcabgFeVkJf
Hm0fPmkMTWNLDDHE60bXeWTJ5XbuiAOhUT3NSJpoBhCwXXDKZRIBFUQCvmJjGDXFTyepZdEw2/F6
wOHAepjkNTasVGs7ioad3M+xu+1gF/Mbj+4uzKCaRkm3IVKFiDwA1gYPBXlcHdb0eqcBhfnfWxoT
Ag/lRWrlLvfI2GdfAf/X3PB4kvDR+sgysFNb5U5p4EnLwbmtYq1GFu+5UgERbcXJUkkCS+iFX+yb
pjF+nqJaw/UVhsx2ZGK90zER1cYBPRfb/TNV8bl34IvsGLE54Kwz5bBBJWJVtjfPomrkQO6Np2cg
98zox5IMc4C7RjmgYbHEMrVJGlCrf96jPCSTt9rZhquhWixzFTFIOno6JdIP5P0kpiGC8kTkI9Wy
sCJ7vGBn4UKmn9krckNDBOW3p636Quv6kN1kGGaz3qiwP8uVJlO0/NEdJBmfB/klCfyR8NH8YpEM
G8XZPBG+4tnKkLiFjYSZ+p5LVUeTzP2BKd/gs+ckYUY9RnKPU2gXb/OHsoC7nzCOmPZTYP+uMd6M
mkIIshGb8nrQFdHHlH5BfPQ0oNA+iwASTvWXzfuVqrYq+RKjbIJmH6s0V2zJl+ZkyIFiouNk3WFm
5Fw9MnY7T3byb8cWX3pljkN/nH0/n9wfVYsr9XWO08vloS4BkEBRyO43a27rfB1AeuDbhDZ21FKU
XCIZSQd57KbZGYCI41Bgh1PT8aeZpp43RWXCElMSLBQZTEIwkQG5+RLGv3DixlyQOxyBxsobfNfu
kota6bT5pn6eHFGyfYUBRjzrObGJrY5Aq38Tc/x/BhiJcXkJQy66iZzL/6RyTkAeVhhP5QEUVC5H
nEGTwT9QZRnQ00eX3cM8T4qaL167bg64Nc3HMJv6NHSLhuHMGsiXvnrrdIvDljT9JhKKeBE2p1ON
VEzwq+iEB/7gRBtP1An08QQOqHlN0SESE00ugjYwy0EB4bsVYRJUd+mapmbAAcIySoPSQ7FBnFWs
cCSloSa+O9FfpI+XUkvOq5mgY0CryaJNjf6xHIwJf6a8lH2M5il/d4+mJGrADcDAVo/lxvEsS04z
7/P+e7Rraa4Rvw8K1w7+dDiXe9qkFPMZzoyP2durvD6kWkwIbkBToPOSgOFjgI2wk492CfEqvzko
cqf0KpoEQ+DCF4zF7sPujpwz/fJlF63nVbjncs1FZgiB+OIB/eT2E9RvCNo67ggbtSiD1JTJUNIg
o9iojp4ARlPdEy7ECOLouTM0rPYkyWHJJHW7vNiNExWkF5HRxItp119ccGLf1E55+4/bhQPCyf9h
anAx9UUvBgffQkMz8XFq+BA4sfE1ACtKGFJjIQVyU9yr3nKrggRCztv7qqsJEwhmpsICoBtDzF0N
mNxqjO+I5HgVBsephM3yFXXxGKOL/Fwklhx7ZbOp1hxyWq3ff05e1TM/ecQG42sXYpWfyI8J5+ON
JGDH8QqqXAaNdIApiS/VKBpXQaCNfq5Ln1uUOy2deSSRo5vOSiWkQ/HNBnVChViUSHMyc5uuNbcx
SZuc86M3IMQLPMChI01bP4ch8BjPspOyTcPJLqRvV69RDg6keO9Be0MfOow0gUIDBC5oOk5L49F9
cSySmYZMTp3KCOSfliNqd15SwUj7Odsw2E+wteWW5+CY3Zp1I0eonGLC70gm8ioZvBGrr2q6aSoD
06WBgzDLee1PCLyu+0Blbz9+5ZdIifpESKz8xSsZB1z9Gum4PH+8uHtX5DSeZdqNzE319K/b/o77
hHRGBca0zvaiCEFTNJPjtJBaMAXBxaDz0i0FDUqfAHgcX3+dEOX6HMxMiSDOU03rJ54P0x9KNRC/
UunaN0RXZtEGpVIUtoKM66lWawOm6Qhccn32p3OuI15Pih4kmFOKV8xNA/PlfQqTK1nZWG+nYvbt
EvPrF0HiV+EvLxXv0qfYeqOkkVea7hYY7SIMYCc3P0O/qV9zEB2dCpVmAs7VdKk81tuVRJVTVqHQ
dv9jitrevj3CslETkCsEZ/sCUwnRmXOpofFf1ncRzgeaEwese4Pxnrwheb2qS2x86JJu6ZOW8E4R
MnIb4ZvYnbivrnsQCCPWXXj8sWaxQfDdcEVzbpsEm24bbHo7r5AwsLkZGC24KcmHWEIdtNzzsoZv
G1W4pK3yxqcGNib/tBcimwaeTNMy7k2z4/BZhjriGdL09bE0vwvkHYJiSqf5FRZXJYwyfbWlY3Cw
9mDWRTFV3OKDIVgSn0GHKK1McMq0W+1iTP2MLk/Dz/h1uGoK03Qr4/4f5OHM8FD1oWVKWZcUm3rs
7RvUB7x2L8RJEqrj4bKoT7RSQDS7iZJTEWgvn6tTX2oq0Fnfsj81WRza6yyR+ytCx251Rk7vSj50
VC06mdCCZXolZkl4mtNnX1ZGM4p5GinFbtrBh7FrWwxqokOU36qtjJRkmjLSm4gC5HrlWLlydJ+X
s1k15OtVFohXqHhu3F0vA8IQ/ydje+Ig6o4RLwWVEFOzfJiSQoOYgAse3LIJ0dD05vfhhKjB5F3K
DqivQdvhXMa5KPC8oyBN+kavz+Dtq/ty/+5asd+F2a2g2zIM+oq0PyatdBNEWpMLwdXh/p9Ttd2I
AMYcRPjLr4dD+WNWdwwxxUuHWWDUEnL5rlKNgKxlO0eLpLMxSM73akAmM+LQhJOhy5YfzLz+LylR
ni5tRHY58AWMC0jb4pweDn8QFAfIqRsaHAIT8Fp9MAkmDoJnP4VIUJ+hAn8P2PXLXPUIhzwyknWw
qlIN9jpz8l83piYeGFJnDJldcyrrva12/s9DNHqxkCkwYZhk0TDhJCbdsc03fWOgbmhr16WLsP1n
RO9iIp+UdrFopCXxWcDcFiRWZ1GwTG6o47B7umKswNW0vm/HguFa0uCIwHhS/hwSKNjIzxAkol26
1k0342p/m/gd21loHKXmWbDVk97fPUeKQSjkd2w5r8DZrXRe19zZVGRGH6ojryYLKwoDyTEuJ/ct
aIqBV9jVREzp3KNC4vv8WTRJZnrBl8NntPRk73C1tUwj3Rf4Ns5nP8h5DXg77L5CJW8/LhOAzB+l
dpvMil1msIZ0YSvdynIsQBMWlQ8+buBjRKiv/kmoNzvK6O5Jj6JaIz9rm4q8l3Sc1gvMuUeUEa+9
XDn+o1loAFpQG2P4mLKMs+7b58UwsCXQbFfg5pX89NVVZz34B210C4ldgbVspoB/44xLhAiVb5N9
iuAUAc5VWz5auZDqTc7jiyXdzYkPi89hBbOVEydRrEmKVy697f5nV4c8JlRJARD1U/rj9qh7Xp0y
KFABSzZCenT/db8qv10uVVDd5chR9fKXXOHG9KsWxcX6oQYBDbIrFJ1WToR/vXjIohqULZioNSJ4
XXzA6pNQFYSmBV97q/6P9vdcH9sWuJxCKWO2JdFaVuTn3rx6u2SF7DN6bSOxUVsHw2skUH7MoevA
KiJsidStV5x8/E4QBzgoKijSQhxxStp6WLDpY5u6/0Y90bbWNhvRPhvhgKsLeHfSQf/uKFw9WrHB
fUFhgsejKl7hOI40DhzCGjUBdTrOl1rzJTunYm/TF3NPHcG203So8/j9M6sf6Hqgg14IgMsKjjYN
kU4LD1+JV/a1aLhBOXUa2Lo4Ppgb4cmkGz71Rwu950hSUWhwtJaYWIMwSrOXCsDdyXOGKEm8Z9Kq
IqKho+dY9GZj1aRAf2kRlCxqG72AewPn/7rd1jSXM1bk0x+GuB90Bpb4rJL2w6aaD7qJWYzgs4Ak
kVyCYMt3eadWWYYN7F72g6v7ZHZkgysIlU8XUBSOsHR1gff+ZuSCGEgYeTqcXdzmKfDir3nJwyTs
lF6KKq7NCKo4v1hzUs0rXn3EpTuJ7K7Bir/iL5WVihRGMcUTfze0NIyv4LplMLuyAmU9WQybQXrJ
bVfIQksaZ63rPEnj2Ac0BPjf3A8QupapYIQ99CgrMMJPjy5S+WwjCdPwEQl/WemKDzcsxovjBViL
L6eWXecD6pTu2+Cwb7wJbgka5MRX3hrQ5J0w2JcVYKwRpBIBszUB86j2D6TAo4tgyS/MWCtPcal8
UV/ZRxm4giVhvbO3ZZPIwGIMl2IpsxAn+oCcUly+Ock6GkJmoAnCN4/pdit8DonCR4kSB7sGyNby
7bL1KmvjTlviH8eos9LxFzGUaGfzLY177jdQbUMjqAcx0C8lpW1J7o4OU8mbBRBa8/3m452jZEVv
QCYrYuza9KtKrv2UxbNcuz0EivYxuBS/bImjkNJGXSRE7a5JqUe3W+u+hhKiObZGYX2eIspRp1Kd
XvsPfj8xfy7kPtgHIDgIwQ4uzN2ip2wudixiSDbrMB0kCPCRs8J9OXrhbDV2cQh9cxFg2WnYMZCN
8TH3UbfN38sPJbLBFbMzeM6Oxs19nD1czoFfiiF++n0PbpV5K8shHMqN4LjEbsB11zcQ0Kdy7vmQ
WPf2f/Cza/ns5EFeqeL1jcaABgtkGXqb0sTFQeBpyqqsfZRcDo5EVWlJ+/BzKgyuE7Co5+raelhb
/Pc6/Q8EatfDsQj0iKNHI9g+QA7DTzyyzKE51oFRk/3ky7WH9fvn5zwPuz3683tMoSld8z7BJJZh
DDqdj5vb/etCB6lOfBS0xDUrwQYPCcRoUDE4Wi5Y+neVGxegJuJbfjIN3giV5FdFQG2C50rdVLEL
E07TI9xOCHFzbK8aIMtR85Iupx7XPZLFa/uZWmDGj2WA9+S9wiriy4/0YmlyNsTMi6z/UdROKnYP
qrRxtTr1KRttKgeV8OihcZG30Bblsms1/00Og0+Fyx6rslkefu0hApzeYROErzMmhPbCPuO6ZAnd
4s0wxneEUnEUicQUQsiAk07CEHrFFUs1UpWNXF/84gBSGdanASwbbonmDCAHV5PrA1syd5MGL+WZ
C9AZjEEku/QnrSurbm6Lp+YDh7VTd2hjnBG//bIlCVglRgMC8cLYHQwzyw8ui6m5lhSvWoBeZajs
cyLnp4n+yOiF0S4LPw4nhLAFI5cn9ISkN0gUJE49nBT4/H3R9NdMuh7cE+Vh7HdE+OHqDqur+jDP
PKP7+BchqiBUXzXCLellpAKrxkBTgCsiyjhrp32AsrlMjNjrqjJL1+DCv3uyQvfQHnlSh6b+1CQW
A9kUd5DXGqfnbUOyfzITMg1IJrDrahSnvMaYLWJaq4OkVo0YSCOwDgM74REPIvTQxp5Fxpm/14qC
SbaDCNjwNn9cD6Oe2z8RnyyssnQ3sTRkybdLRfC8qdqqUwvQgZciQ89Bsxs1Fn4LW6MyUWIlmOyq
3NkSVw0CDmKIxdB2g9b2wzoW+2r0fwLecsVrNaNw2aAnMFDUPiUEojv7BuCxYZa+IC5Ow+A7iA0h
3laptWLMs2t+HOSIsYecghJOi+5MOMou410+XhwJqaad2eLhXpFZsoOVhSuC5oXY6PA3rlOdpm8I
45n5kd08EKeXm1clDWuW3K2aWAfG6+3X/cyhRALZlEgMW019xMFmffDRPvK0ZnyGYDxzrN4z6iqT
VuDTHVL0s7JmGA6QeRh6qKeolCtCJ9CkRnlF1rq9x28myxsm+7o993VHGrRRMN28+WJXeU4vSVvv
+QDv4Li7PuciTU5DMyqpTHz67cLBUvZOHh8htX54e0cL74BPMYyMKk4Rhp9htloB6858h9jrR+Px
kmd2fb4kySxmm+8L6kD7iItVqo+MB6SnB/JoPnVwdWm3YVlj1vHrMh5lZjnkJKkSe4G+ncpnUAwe
PZ18YLRrp6XQnRk03P8eEW/RB6xBQvSV79KB1uw4zgknsKgQEJFZc5glWwjDKOSMzgf/3LXDS2z6
f/b3sMa2huIGPrUurc506O40KvHo6oKTxabCaRB2VsAXHs8zHfmoFMhQVXqH4FFVrFaENKmSYQ50
5uDUpy1ThOxwjfkXy4eDoVi+ngYwo2fltiv4SvqCnF/cp+0PyFAqVCyb98r5PzuwgzurkY+zwspA
eNvo6n5B9p6L1SYx21PrxEMem/yaiV/YTt+bFnWZh74Op4tWTmjFDe9wN90X0a6f6UJkaSBMWkZ4
JmyRzb/mxc6d7EOxE6AsrQCeeUVouyvP2DbcVVxwk8D064ANe3ucGJ4elCsXno6+E6jDrRkeczsM
sI9SkIJZwBwRJ0dqhKfcMkB5igRCO06AcDhIoi7GR84Hrs3UGwUb16Ms2IOc0PIYAGNY1yUqXDkY
oUXvRY6AHlDU4vr4M9+8Z8Q+hq5V/9FgbWyys4EYqXZAkStPp7SnLOmdn+1DxIJtlD9DpcFSWqJ+
54DlDtoU3vnL8nmNYTk4oe2KK0deFDTtmm7hJXCFG6SRdY6EKAUcKbTzf/GGFmfqu6Lr8/TxkL/U
Fy6VsKzSyDPWCGsf6111y893QHHG0mLDkM5JcigsidVAf9hcs/jU/3FNTQjRPP6ySBQWDT3kV7z/
KWnnh7HzyUo2huNvds49R/zu9qGnGQrDHcBRJzXTHoNrAjU1G4uTTFt7ftioTtrSq0mpIXixGafu
hykgeJaskqArIXCJ4y1kpoGmSp2ffg8fvPIXtxL+wSHMk03ljCnPt31ohAIvNicMpJQpVeP2k23c
16b7jbbVI7+sEKN9aYsAIIyfLZqQLmtUHufbEh9U4sYbDBkgTjAZo7DWJN0SIB7zwMUmJ0kg0S1i
Yots3ZIvnqxCOu6huQcHNQG4oXfKqqJZ99qJJYdZSNpQnlAWwT3s5ZCfPONFW180Xcn6+9iLDx8U
pHBS3cC8VgaFOFtTGZm3+lDZRnPrQ7Gpufa3CuokHBPlg5P9eLyZPa6o7t9P7I2Aa+8KKFVzNvDN
wLIhYtzjLXLvZHVYtQx4l/ujDuDFOtHFAMPfVi5uPkQuT4Vix9ZFwRhltOZDmay5CnScCm9gTpUn
075Q1+NvwuRiwPHC0Go20avdrKsMH8Owe151UGbhBY5UjbhATUQ++lSQYYiSTIjvGPSrvxAOIOul
67eKKnL7iet6VuZ/wCnGD0V7tpCp5jZSzqvLYPDAIj69or7HTFw0eog265jjAWXPCfL+eUf3TleL
LgVCpRO5nG3DMGUqjF9mbdpuOr/GTi0YfnI6UZImwWDcqZq5vZHMU8VMIGb50oKJBxmpNUxpdkIt
qPtovIIBf2KC1NVeG1fcw98DCo3khOwZa9SsDPWJAIft8MxcJtQQn/bSBCnN4skoti9mdRhlDvKa
XAh+dQxFxs/Dt/H/8e9moVa14ir9eQDw3VF489o/QXkUHN0bZ7r8vjedXsbrwLC2sZ5DerXdj22A
y7rDB3qIMK3lVQJBZkJZOBbOHdYow1ZJt+bbPHZGXPhWBy6KbRmUOZ9OFyi7UistJfY7huUIf/si
GPKEpVW24TuwrkbOsekZF/SlLvPXk+ykJfcVrVJFFKmDdEuqpn7uOyrFDB1im4Ib3peKFnf0LA7A
TY6RYAary2C8jUx7cM5bvg4WJlivzBo3n9GiwdLIFzFM6TzGRhL0glKDqnxeRsrvcUdLwOYkEOsw
zvOA4iPFKGRb02CIp0bq7lzRQQuKwo42RtLRdcksIoW45hLtd1E6o1V4BSHaLbV3lGTu5j9djXf2
blndOD4j8CDXyTc03rwnrbS+jXwLl2wCNSy2XyIgVOVR2ZkZC9tVcoENiE8Q+6qY0zmLL4OSzFfM
lsvb9Fral9cQISH6TXBoPnu2U07+fB4qa24lacHwvqBT0VcOk5bP/uXJNNrUuYQ9jWRy5vPTFZqp
TAf7hwNoqcTiyyaQRUPSp1F7XtdI1R2KkcwrKZqBd3SwDSacyMo+LGXCSXpTvXbIW/DT/YlM6vRb
2hJ3dSNzKfD4hVuKMhv+TBrCyLiodp6DyM+WYdyZ5eI8F5np2H0qjX+DkMIW2B4SIsILZdlYcvv/
WlqLet6mqnHFtgdpRMmz4QqsB+S3/mibmblM4otMHB1EDyVpOHFIWBypmJfwo4hTywRC7leXLAA+
c1c6m917pCvVLSxsRPMgQBJoXTDBNoIGNdsptMeNsUFVSt6YeuDYEJ5uRtICFMr976FoTPWA21YU
6KeL9KRpkQOllfrdw0ljGDiOq3SoLMlpy5MXjcFGQjFlZ8d4N/2qkakT6HvWfgyy31fwrCwBDstQ
flMcp80EC8cG3p/g59vQnTLklm9svrHUILOrFnEgKvYFUZ3CazReiTitaS2tIQfSNk20aC5USpgQ
YJktM6dX4hcvEBMZ7nidoNpj0ErtYgGGAhIwHJCjfunGR4WCIH/RX5OuIs/PqZANEZmpx9mwSFSd
QDMBxy0d6zuncWS4/kbzIkg68ImIh/RqagZKParT/p1tGXDpE//pCqK/Wv8nw/qBTPZHTuCb1OKj
u94MxnF65jagR2gCoh6OkwjsUi8dVIB38zAX9mzN/cK+A0OM0LCgYSRZAShIEPjT+1Qmu74QeyGL
UYJCTw3cX7HECgVP75LCWwqTywFt8RURY10RiPWKAFGH3kUrE9gJa0wmx3duvOBYsoMDwLNw+N3T
RmwZDfnh3bhzMqtEDepRUksvmzdLzUh8zOjusWqQU9vEqtpzZj1bRDmAFPgXCrybMQCnG3z3oXHG
e+Ya/6NbKJj4Ui4EyZD2eLbhuR9F+mC0Q+FuBUB7/SywG24oGRwemOaTf3CCxvbq7GN4pnwNjuCV
+jwgqrXDXSrygVUI9CejoRt5uz7z17W0a3clBNquL0PxEyiJ5kAdz98QAx4pewxoYYAW9KSNyJnT
CXB+mGWOX5jdKkL4jNw9Lod5cCCZFV7Sk3lHlo+B1LtaNXZu9UKbVO4HzPGvVASvDtDHCko6RgiV
zmGTKOHkr4cAhCDkyeYyGq+23ZmT8rjL1VGUghhv4pQu/9ZH5/YMDLh2xnyK5URa1LiBCGhNCUTv
/3wX78spjZqRRkI3+nfQeCgjw6Sxj44by6jcBRcZcSudPOYk5CsSsswba9Jg4mKuEIXkjVtSxfh0
5493XOi8beI2B0230A665m0HsJFBzA5he5aNs6rxFKrMgC+0Ubti4FMm0QLiibX+ma6rIEOcbDXq
SyQsg8nvxdIL5vNonoymNVQt3hJiquHdigjn5Re/ptJDVqbjzmr5YN34OLc53DJJw4kvmyEd05B4
HNqoC81tBmb0pYdZSKG8Ofv2W4OrEmtBln3BvWxmbZPPU6x9NywhchPIWTbd0eTSZ+Gvz/6yJ06m
nQAYffESFm93Zavp4dJCyl/9GkzQ9xIc0yN1h621DfghSGvEB7Uds1fFZWnkgtk5cII2vtTcHKwf
koJB3onremr6QVITJ36YAD+ih0spQOrutDgmxbXPJ0BRo8YaghR/xFUjZmF+6cQMBwlMkb5uQurm
T+vNsF4qkRCHSrnZqLka7IrAfGCMxmYEpcI7JGmJ6Wk1z0GtGfxfb6nf/ct73zre5kBU3bHX1tVl
4/rXUqslRQBFXogfu9gofjcvRDCdWPcJQ+Jpd4W/xYhlUnJmvMtGfyOpiHcJdpZ0J3l/20Znvv2A
gxXsInYtnKmMYNBD4RSTazYwK/K37WCawlYwDDEJnJ6t1fc5U/UdJ6vGwd3WijgWXn2ko3kHSVdJ
NqleO1qslQTW2n3cONFKoercwNyQtZ8tDtJIogNbsA6NdJOmwVrxTpDNhi8Lv8+JMUw2RJzL0Lqh
PqvP/Nkh3ZLO5GRgKRIol314aNvI9Df3lBmH9fPYIH7WswLGKxhPbcPQoM0a65BpcUfKjU6H1Kj4
vFsR0Z6qQJ1JBIetNaiQzYQzyCK/Q0PPMNJmOMP8lHsXBLHG3uwHNX0JRo7TlBpqbr/a2pXco2+5
n28pRwIyLzK/PK7BsDEHh5gFOC5GRaDl/esmDuA0bhQD8B3+QQGvJ7OHvU1bHVo9+wDVkW8l6lBC
wfg+XHeR+3UHdWgEWm+ji0YKzSnUug8QCYxkcdQoYjZLQNWBhpNw60Jqz+zNX+86gMhjNjlBVJPe
2mqb4KuhEhj51VKpL2GHen3mmYhtV/9Vb4YECQEa+PKQ+EnfiGosaU1AV58456E8XUgdB2f8dM4T
fShLDngSa/xPeXOjzMnXv+zyaG7hoaasC4jkC4vg7h71r/joJ1QxIPovj3LMQFivhsg0gTYEYzYG
C7b3I1J2wiFtahy1iOMGrwvP+7H51JJKfea63R+Yp/cQM5sgPLA+r+Nx7gHIQ4GVbDKotc9F7S3M
F5/7InyxhuBOptjyc4kfWApFlT+RAe9mNDlek1AW/sIvRMmNErwjBPHBVdvvKBgdwjcQIJ9R0Q0B
hx7VFEs2cJoYROqvQsxCE37/urogTV4SsMOxfUz2MjxTd4fYGiiLVq3fYHEuJnCPhL5yYzid7lQH
LNJqK9CBJ/Bai2HsYxIhni0cfWGoAh89pQvrB0xhQGIaJ+IB61LSCty8V1sTW2HPnpc4Un7TZiXr
ggosb9Li4LbpUE1835uVWF+8uDsBhevvzenDq6F1d8i7PjgWmmuH6WiH4H+Yr+KTH6qU+mOOw48J
hHLnhhKRLNPONCBky0jid63nbyoa/rWOfp79dpQK+G89/u5og5owx27o26Fn0TczOobPsM4nMC0Y
x5zxQSvspf5AxXHgCgTVe6tfWX0atUFats7W3tojHEwf/7raMwexduGpH3RDt1oi1jyTt3ldcoNp
8aWPmevd5Xg9KLwH0MHkwuf5pLDY5UFnWwKgWwtYF+2h0Uh2V1i/Bfth6zTqBEAkg93idrEFfn2q
+vwaqkoK/wAIWd61oujgm3kzq9bjThEOZD1UwJn8Ztw1r94dm5RDs5Ydi/oZh4nTJGSMyjNvN/Pk
Bwpzuea2JOxYsQSmSCkyEAKzJrg7KGofDlKdCtDUTw9Mylu7xv6f7AY2YPp1oDgpKpzSkaLBYDpE
XZbqg1barooXGAcQsGD7D75IzzJEpt1BkX1yOqCVx+9dCIkGHajFMxQHFXcqk0UAnn6MH+AxFl8L
W2Qb90Q5LExQ047GaGqsFej1eQAXe3EiatBo+nSeQChsJcgplw0vaWHabdswoqRKXiBvgZsPwpTj
zZlM9dDTGuzybrC8jrtTk87+kGA1E6ywbHUWbBdXhc5/UaHq7CZRfocQzer2CweVy934X8sQECgw
0TaeisfNWazo72cEg+AWJ8E5dsepMt1JKzvuEzyUX90wSAur941Zuekf0XeCxPoDwYXUKGvj+HGv
VjCZb3u2R9JmisD1FuL+CsQpiFIw6O471DwOLGoTxzVkI5467P3yGMRseUZ4+Ykcolvj4T+0PLpG
UCiwEwqslO7NFxEnJAFpXwJlJlYyUKwL0dhPcPKIxC0Fhwjm8QWnk6neprgBSrlUXZhin3/aGQbQ
bMv4z6FINz7q9nqXsOV6k6r1z2PtEzRgekzvq/BQbEF8Gprk242UuoIev6yzDUSsR5hAoI+6IGUg
SX+8x1dkaxqtJr7c6aJoLbmRIUuhAsHC3/twiC3v8hihgwE5P/M2jTDYErmW3wJzI69TMQvsTg0w
TueJEFGf7jbLUPJhUioYGFgt+NF/LVwHvn/mKMmcl1voSjQgHlcLvEIbCLIXr0nVf/oyxeNSMV2X
NwARSKOLxrMkRTm+0MRmRvcxicki+eeMurE9E3KlwDm5CS+H6AqORo9TKK+CZmXVmKzcCCqeWH8V
qmFw1RJ+g8PuyIOflfP++Z2tohnB101vMVNwuXusQJJvYLLyPfZVtVbjzvR15Pp6RdmcyCu0i5K2
l6isBA4/5oKKfScyyHhMFEy4MjyMngMdOoGyIz9S7pIMJVOr25xQUjPavGpfS4aAXtt5S0snw6K6
Z6i+Tm+rvNfbTFcoQwPaumhbdwNHqFV9d4emMMbilhAxTohovympSTnBOczN44OE/3EQ79r8H3Y/
8wFXGxjnbFHu3ltJDdEwNdEl7EVoxDyMFtIXOezbpWAsT8EgYa6eJx7/JmmeDl5RbSJhQkwc+NJM
oVc4m0ofn/yEzTI1cBeNUjQ0pEs+rJo5/1VAviuRxdIu4/g99bjUT1qJcFTbems7UFPCKJPHkxY/
B6rjjZMMrIb4EtX7GhRJh+i8GcXtbBp7Aw+hC80XRhN1FFSUKz1guprJ+/8+v1H7Jc14BwqsGjQc
QhpkOAIdS3/FN+W/ccdW3V337UXFxZw0/DAhy/HxWiDK7j9wS6+Y/BRuxqowCiIOrDtWrmRwMz13
EMrIeiogWdA+2G0Aaj/ED6jMJim+skUyNf5aMbiD7zg1jlJbFt2Nv0N+Q5jZz97qM9Jv/Vu/zfzm
yY/PvOgndAXq1/J3xhq66ynIxiNMMPC5BiANJiufQRdEjCwrCvxqniuduHpeBs5L7ohd0PkAv30E
u6dZA4IRpNx9EgvQhLkqzcHnM5zG+PGWDelu3WAN85dAD9uju/eifFYnoRIcxzB+Ye9RbLMul8zI
5ePUmycK3404wtAN17KFLEdxtBg2qxfGyJl0bcct1Ha9UlHmpP/Bw3DslbBBPBI86zNMzhHZZUfl
kd3+M+YVKZj1aI74RkKpVD2XxiPFGbAY5wbfqKsx7bJ/RE24Ixj5H0E0muqgY/xhQI64dmTQCY5A
mLFNKxqfoUGND9L0ou5K34+EgwBuCdsk8YZgzB6JBO+aYhrtdPPGGXexJDsPZG8xFWjj4OjGCI1T
qlz5UHsSTCYK9fKBYDRrqZqz7BTtDWpcsRkiBCilJ1ZsE8GB3FxT6+1gzCvPquo1m8Y7rjnLCNyP
44b8i8b6MVvMinomv21y6B9EdY73S5jKIt7hnJqlvCOcKAJWOIbe6DbSGkoobtfTVDJb1cZtgXGR
ugJ5OH+d8k06PdiQULX+n17pbdTQIPCX78584YRWr4mD5KW8mDG+gKN1T8Gh9nzUEcCBCPzmGqpl
m9vJdmWgY46QtDOqmJhYtt6AoUnrFL/wnLcyq2k8abp+SLOUyp5NIIVouOr/WUQQlu90LiE0Pi7W
OC6J7XCGl//esonM4OHO5zSFDJam9tluhnSKwmH2AWKyBlNhBa/N5Sfv5L0Gd6ndmT7HZCJrhRIB
jGCrqIbv2/x1+C/pPqmXsHwrMJ9M1uC3NuYUSGj+KQt7j6yVsOo2DMeq9HJewaYFjd2t/bJ4iQc3
LuT4v+2oBTB1n/SU+MRQIHBQHa6IJlBxMMoF05Ry7tK2OttV1QtPbRgbl8TTHW7IOqAvRaepbE2d
CIj60r0h3lBDTX1G8xj6GXrRhFi8KVuAa6EbbRj/xURc60sQYS+00JXLPNAN1t6hXo/tVhbxJWgJ
0lS086Nf1w2tFtWMdCd4+/2YWAwezim4QCWFpI/5QHkdRmaG0pBr8YKOF83v9HmlNkSLKkW+o8RP
NZUjOdKKEUvrXaOfgH6WvQI/aZ6yMS2PDDBoGh5UkIYYYpFxaAkngGHl0lwLq0C+ptJI6Knj0Yxd
/WzDGMM4aIM04dZRsEzEWeSvzIG7PPYV0re4VtgDh8B6Mq+QFGew8BXMV5YPcFtNi9+OwOwFO3zT
cmQOQfuqyAWw70m1jSeoZTKCKkQy0Y/W1WNGWjs2ptEGlURkygG1W2WSk4SZLISJe1klZPPRBcFf
l+yv99noDXsaFD+t50CbiLOcn837Y2xwzM44ToIJ01sXSIePV6zk0Oqec7EKC2S4Q78ECjs7+5Y5
TpDnRc+FjqDHQZ6x4beuOXVoL2yX3QXlqbp3XMltHM+ruj/UgdT8Or2OHGiZUu44HSwzeS36HZnf
po6X7eb00KWegkm8AP9c1b1EQUBdQZZrIpQ6tQegWn8qmwPZ0wikJyLpLosCAawnaVqe6uoNk9dP
AR1gvCtRhsw6IaFQdJaa6uzaG+bJwgou2mpcNC3g0TucpXnVtm/9VcsmAr0t+PSAjqa22QqUqyWO
BPbRff6X3Vb57ObO1V5rlW8Bw+tu6ncX6jpPaKbDCZ6QLrHXqo6JaLJRaVqpmmXK/d5Qlp+ikmye
YAl97SIvjKtJ008j3g/mIhND8tzIwo4L6MjDacTA1Qbkg33kR6wrG+tkdcG6lVOMJcqdlRE5SL/n
naW/iNq3GisaCVXZdR+Zz3drgq0a+td2LTmmqiFcIlqgHuCINY/Qcg/PrD0sAREbt1eI9KEZSQX+
Auc+9OVSf9FfFOGnJzwbwWIa9smsGcNE/mLlAME6Pv5DBNUx7tm/UXpvv1H06LT66QOKDd7e0L0R
rjo3m46qToRtqHEzW3th2TbmBI5wEdOlRP6vJWO0p25ZS4XZZk2JFus1ypdt1zz0zaiJIfMuNNkV
w06Rg2z6ChZE8kYrr/EQBjzS9FN0Z9lm6S9C2YY++p3KxNnks7ztSQcuUWsgLA6cMqTcRAJI/rrW
zbP79NxrcUYCQ5ThiSBtgRdFowEAB0y08WY1bNU4QBIsA50YDjX3UaDwez8wWon7OB7ld/Va6r8T
d+7DXjOs/yH/S8ooNe+y+eNfc5oHfeKkeosgMn80CYABY4o3qIPABpqpw2uaLYvxS/NPbrQjkZlV
uSuWlp8vG5uXNnXYKKPi+xNjVDIpfZK2fB5I372n4zftLTYXtGgKhp9YHal0/Yz2pIpPbGSt+D1a
2mhF5z1l6xmPLPm2P2H5QrX4jey4hrEubUXNN0DGmaeuZjL4mAYGvtw6z4oq6QqvUxv/nrer3rm/
BHe5OaAlGcYPxZpSwPnVouI3J3HPkrPt9e88OVyahIoeWc6+SukA050ddwCGcQIiWVcnJe3+tGeB
ii03zFBX/JY5B53gFKYke0ecxkvIquLcObgkALCTr8dIgRJt+Ys+gBxtQUrAzkFmnd0aj8F43Oic
DhrqkXY/NxtcBrwjD0FVZxi4AD1yuyliH7r5UGPNZ4SjHWwMa/T6B0XgRr9wYF5dLe0vVTPAzmNn
hDTN91MheQjYvpdNSgjjtuYwjGVkCOD1f37vqbhy+UYoHznFvtberoHOgzqFAxN6hpfKdXXfYKWi
azq03ZeQdKiWJQRaoeO82j/OprMjYZdxNz0iEARxBOMWi8fZ/ckU5pR+ejetLA55vU0kYChqKi3H
CdEA/G52HWiE7PDHviIedpWqE6he/u6ywLHBWEtmtnmtiEp7ENViqWSnRFR9fByex1owGtWEX6aN
obniqSCimPciffvNQPgcBEPZTP5RQxVWCBHuiYxVwokxvh7/Bd+3bfgavVMBJTHjjM0psoymnuws
sa/rt7OVHfAlh82MqPd5ODob9hbmIh50td9OjaIS8ETm6kO8+Fg78u1vBNUvymvqNnQ4FAtelli/
AK3z9JEOnR+nvdTNzGERBXSMfbnVjWzsyFQTrfHZUD4pQHbIZT9SRE8luMRH/y1c+HH1h5S7Y8sE
mNS6U9UhuVnD6zcSYrx1GaarNBNjFdERGjMoZaJHH1IZBrZqjATM3K2OlDepESN3P1NNxpsRTmP8
EneUpAxRY9UO1BCI08A2AE1PBns6Dd4ABaW6fZxnhk6exCh8WQ6IbPqdWbkgh9Skb0acDslKFGU+
oG+vHNj0bY6ua26pLYTi8odUPk2D8y8NMACtkd+TuT/VmjB8dk8C24ARRmTmM1z+ykbJwh4AlgAE
LS/jmwXfMYevhbr1E485RTaaMzh+YXUTj2LvKmKu3mKCSkpyskZ1kWw3010HkY8rXbHxlk6dy1DM
oQbqzPZjarvJ7ad47QmCDncok+zlbKid6AI2Kih7hZ817vBoL9fijVO2rPMt9mLcUGT9+AH2MWLk
UYkNV3T7dcU3WEiKy1RmvTFJ1J0qHaMIr1I9oAAVGvE4r2iBnUWIqjmfUnQdLBHIEgV4zX35sHxy
gU1ljDdAxf6X+j7asNdTZHI0QwdroALcaSEeOSPXIC0QGN5A5J5UyJ+CxRgaDsmS5k8RrSN8lwZX
zeRhDSu9Luv7qn1Mr3WrwM/6AQLtWfWVRjYKn8eniGXpvKWiU1VlVF5oh+ZSVKRf/qfDNIekCIS2
8189Ba2/Xw/m2d/E/zKcHM9fEC+qTPkZETmBJAfwRbegyrUJBzq3zveAvmdnXyh+hCyGR3ikuAU7
yJuNNhbGFIJP94v9ymtatTjCYywTwpidTtXRbkarhGbMnLTEJTsrZa9WiWdOnmbcX13c2OoR+xgL
moNqUrbjvugYseEEPkc14TqvCr4bEP/jlxio6XQDcft/wT4GRWNaeollkjoCvPOupcP3YbwL5jBJ
pa8fDx3eGKW9zvASR5m2Y5lrEIOuiBAbGuQrsqSAcNAmpJMwB8GaCO5wB9RCRZ0dZumTJ+uUe8X4
MjS3VDgyxLsdhXA8z7s2y+gWIqVKnoKZr6rfwuYel8TwIStn+WisNT+/urSj7ZWlSDXKX42NpACw
hRpxAotqKtlre2tHj/6o1ALo9WJpnyx4Lugam70JT+DL2Wl8CgM2YOYxi7CwlucS3b7FPKJkC7s2
uT0PW8WFbqBqLsAqUskqyh8o94kvjOXlBOlZOs6JMKpL8oHFebSC4Qww6WRky8CG2UR6j1e+VtIF
9iMf1QTPrh2mgezsaEXmB/FOJ3ia2RpoVz8ufvstUema63zr8uk+2SEjWnLpPDgzi4SPyTVgIHg5
uoEwC5+LquMxEIWoXr0FSgV6SB9GTeNRHUPr1ROI+edjmw6g5h6+3OYk4Pm10qrs6ZQaCBiVvhyE
QdPwz9yUG0StJStrSZuki1fDDhy/NsFBhi+Z0qF5rSiO2IQDrHmCL6ZP8FlFsi8+2JIIp7n4kYqp
kDJafNiZRu/20zcT0LJgtGYgY9r3UsK7bdiL0SXnx1la8HUX2ZXmj/Gl1v9vGQTDyi8ig7ta81PM
tFilr71ONPECaRDvrlkomypCpCU8In/KOeRdLCGkjerh/royuyFfP+khtsVo4vS+kGbxKO1hv9yX
iQpagVnGnxIaxHXsmUUmLMH+eG+nrMbz1lcy1n3NyGpbq/GOeiSo9daEQ9a/2hBD0I5Xdiu8dHve
Xf8Geohoy70WgW7xyf5PiJeZwgb3gPKQgDSW7VnvQ+tsQA1yQZhiygxVa0ViIYbDzEouczfmICMx
sSse4iETkrhtvHLfNTWui5PoH1xOc3Ml9Tm4pxfUCHQXSdls5XDYxY6QTSIjgfGxxe90md9b1hPN
HfCetG5ICkLM+zw6xWGVnuJEL8v8J9xr0HDjfUeHv22ssrBHbHB1kROJ9WP+Ks5wAA4KSnDBmQ0+
RcC/IZYs9UyES2qu6yQmjwVAb9dVnnoFnMzHPQ5UZrgXvIyI/+8iZgBoJc8Jpzk06k3XLUAztbLp
dMMtAJonIFD4Q19Lw7rLH+9e7P4yzrWowsIrVJ2bXSd2jBa638v90nImolgsYNTiOpuzZzZ89Koa
GIbCIGefYA37h83OyDt04iOTA+hY2MNoqvxoLYQhBCkOWIXznOuATwrxYl2LtRQnRj90siCSug4h
sCIs9YIxW37rgFXQWnU/nuUu8ZmSueqZYtrFDVPYbO5h+E2FAJdpoEtg7zjzSlNOJourmQpXCW6y
D5OaMR7i49hZhhu0aTNNr9Ff06rB6yyGstFcCSy2sTPpbgAYe+jSNiJdNxh4aFJUg0BV7GQ6XTdP
PC1CBiiRCfVOCLpmG4G5jY3NAte/ideTr7DZbwT26ZzAWNIC+9C+ZgDCW4kKQzTzH+KOpKuJcOPl
oZ2DMaBumHGDGFEgZALh+9M5cI5u6FAsOTaE6y2qp2sP8c5zRzU0s7KuOlD1d9PXetTLczKEjbzi
pfmyEYhA2ws2q5s3Gzz6ZuNdvILFozzAGcwxTrpZKkIuyhSB+RPB2K4P1b4cllDES+cfgxSODEQ8
ihGF+Y+rEuhhNnOYXQicmVCQkMbtBYNBxtHXi2rf/Qs2Uv1w5cWs1Au3OoNp184cUK+uwT8VhwFF
dTUJdeIkbk2j04FqFeLBnPg2pIYuxlOYeH1uNXQrssrazo3z/qnI5fy0qDHTYvsCECtHWui3zhFv
IGxyyfXpxi6Bnc05DXWlBCkV527sLv33BWvqSBEzMq603AVVpCs4D5mjK2fOazmcyW4cbIxMzt9x
wyqEez/Jra2o0A6xNBFmJIyHIFWFiZrWfZm02yu+fcPe2bCkrk8+7dHnsN5IJYZxbbM2xarGvBQd
4NGcNZEs4sbI2fhW5wPqb4E6/7UJyeI4p2CBJDejzhQu3GI6ztSgr3JzXQMm47K6amv0ek7qLhFb
GsrNP6sO5JC4gz8gzDt5527tCXUdogZ3lYiwyHTmv6Q8qTiQm0W2Apvx+H8s0O1VP5ZPug1LDRVr
1EBWMFbycPsPdqUjCW+3FP5qN7t+BRwH7jCVT4rgENrcR25VxqscOLveONODPwr7/D8uutcVjFEL
CHrFzoWCNd08jN9sSgzUvGJ9364NruIXDCLeiZ00Q5OrI8HjfpCcqPyeYV6t9lOgj1OpKBb9t3VB
mzb26Z9WSjKyVfJTTXEr6fIAmMdXRmkvC1SmqveVfAZPk+sdzEzkP7n7KdmFkiG/eS7bwNdHrm6S
WFcPIqS3zKbSR09hlm4SmqaH1KXlJEcsXvwkx/NGv5nfY8osa21DDlvQzLW/udzhWA9cQC6XzZGS
DQLhJfQb9S0IdnEEHm5ZveIlVnR+3EjA+DbpMmXCgO3CGpFbKJShDvY7NQzf5b1PivePLJCc0exd
kXCsBUxLnJ37PHwDLE3ImoHNY5KmRaCm5QUb0E3ysIHDy7vZAWwSj7rSHNWk8LlF9tDukzNmjpTC
Yqc7gnH8bog+XIxd+1wjdfqp9wMAZN0F4cJPZIPMT/QIhaqVjYg2HlThzSXSGJM+NKDaWe/5Ke1o
nR3RoPFfZKEm7AhxcvrnPnFuqlRJno/tJMljDckFLn/DXHA0D5LtcJlhRMdmEWrMyA/wxu5rG70T
YbMYJhTdlAxmpguEqBOs972xn+g69J/mqIp+Hge6nn2mQzcNgzk34nik6SMaWMdYBUs3VTYSPqm4
U+tmw3Uf69KPTvo2TzRukKI40N6NoeIO3Z7jesebDuuXhL/dTBeYodXfSQ1SgLRuT6ceSf1R8pER
FUX09LvzL1gsSn+tw3xqtMhyaz14lTvs7LCnPAuhdojpP2l4+vPchBf7qAIMzLbtn2peD0ByzCoH
PDfL/bg7NCGbANSVRnW3xKB5rAvGAGH+SMhRnAKE4tnGK9yyNP8p6WBzvwfHCU0Msp9bJatC4OPe
nobAcUdAmWBTsKW74eftbfZaLhGQmWaOON+z2aipLW8iLmECZAEKB0vUzjO6xdBYU1H4GCUgHU7w
i2DvmWFGPYd1MWjnvBzetupJAO7X92GzuM4j1C+60D8kTKkQnsDe0ebcOKAE1Mw/r3fqGlwgPCa9
8R1Aj6S1KuiXhPxx8wkoNkj6csWMiS8ofUNEUDhGpB+zaOVFY5goQcWG+uKhvqdrYfIXzuZczS9U
9yTSgmTeZ1PmsUYDypr++i4KKecE+NgW9eQoDJUmHEG6N16s1DSBgXlKsgFyZ0a6TynalYVIeaHy
mRWKxbzVlFS51+/N4ViTzRCX2R+WC9QIZS903xeElM/6QkRFfDYo/U0mVItacLaHBpYDn/CsCmtF
4x4+o4e4n8SR5k+2qvdFPgJQIsFYU+K0J0k/LtU9gigjBP0IyP64EsGQQlCRkAC+SE7i5v/fS0Bk
oWckiFM2jeCgEE7BlwIFyoYW1sA7LfdEauqB8A/AxlnczvbYP9M/OG+D/opvc5UU8CLjIm+Lf18K
Px425kWtwJzuzI8S0BF0XEDVX5IlrebYBDou9dSxZKXYbQGKQeT2YoFIa5vuPUIEHL5FotxruRU2
o1fuFCbWVigCVpfKGZwiEiC+ulPsOoVqmYJa7lHX48YZzo+qazxyzjIaRu5rAFnFa1C/DdzCMurG
jpJkwcsuxexDJYPxSNrVNC2o0ipEDA3mSFIW8Bha0OqELrXhzr0xoSKeyabuLFOZ9oygmMoQkRSj
hTHk6E83G91Kg1nT+Ljli5hXChnU5VRJMBRWhJkN2dh38J9BtQ08lHS5lM80UIQb23IQREq6vunk
VdFrTy8lVoE+BKaIajuYJ2Pnp5TYfmqIlQXS4aJrkn8pKVNhMF0m3UqGIhePxbMENNM93VWYaTGs
Xz2NaJjDipSxm11rv9PqDq1BRdUisIE7ehNYJXbyqJz+pmUPdj4U1PK5FB628iO5stUmRiCIYLLY
Sf9YU/fgdnGx3ByCwZzaoA6IaYbOUzBEo3NzsJqb2apW95XEzMESrslazaWpz9gCjifiqAGwKatM
OoQXZfb2dabXksixUIvxh2ayFAm539zmM5pB/1XlWe7lo236DQ9zPY/VDqfhvCaNBkKPb0FDz1+j
KSVmdZtV1njsStZkMk7QYHqw4NsSM2FMVX+eavoRhgJihPaStP24d4hLGtm9quh1gcDuj0ZQCFQO
lLgjg9Rqb4aBHkQlHmNyeIcsfT0YYk8oSW0u5/noEGzzpX1+jfaBPK2YDHwtU47x2R8qpmmQRrA/
iIVsOtNIMUNDzK0JRpNqgVzLHwpeO93aqtCL4VENrYt4/SUFuX+xb3vTn05mbLIFYQDgS8kLmt0T
Mydetwp4IpY8FtokaHSYwgobDz1SfXBjO04frq8rnc3dIRkcHRyazf4zXLvSyOnBL2G9GwsuIRUq
UVqojiVk6TlqlsdgcrNWsg8OHedUjURXgZ8yJEkxczYLdFCGKnX3U7qwos4ke60XvJGiDVFnR1wx
bPvWjU7QEGipY9xSzDC8XSv0j9V5nU/PcfmcmYNgJGna2UiK+ktUWLoW9V7BS7kvwms2K1SJ8l2y
rjhCuBeK6rm2SmO1RqwuSVnLjXzwzYZg/OmfF1y1d89k44OK8flNpmPPo7IUIPotNPI2+VJRuF5d
d8YAU2AhsVLz/hOiFq58vx2QzPMxwdhOM8y464Uqtx+kNvK3qmOQ6iNsyjpNQ7yl0PHNVhCrdr1k
NBS7nSzC/+CZVWXlXvbWZScQQfrDbS5CBI15n1D3NdNWPvXoRe4bapcrorPRpsWK6yCrvSMm0JrZ
Aq0uC4sJlDtFnUzScwXht1aKw0iQYF+J+Q4Kbzng44Z18jya073A2MZD6nKOWYZ0pyewE1EVipYq
qax6KJ7r2bHqTMKubtm0miO0H/Ee/d6ZJxdYC90kReSt4Av+GnPS1L9GJNlD/zBdblee1K4WUgUH
hFyewrsgFbgRoz1HkgqaBMoWTWl8OIVSAoOEQPB3qefG14+rTjRD0u+b21yQIFwv22wTmBVpN+7H
0A50ORs+1e7ebML2P1AleCoqj09kaWiFh/o6lxvKDleip9vTupmol/kxg54TQNvCept6Je5PKaBP
AEEMpg5HAEdumlrekhiqIQuNfTjOIUfMl61zb5tcjau3HGoBP0lf3KoURcrRsCxJNcqzjuOp7X/j
8huEwuiVR7XdwEw6/gWhgrMtBvXi0Fzt+ySF4F6rcaWqS/aCClsjifSQBy6gH/DDEkYGuhqRgT3x
EJO5X0PjFlp2ra9vASxxBon86P0loB1eYns1K3waEo4NZt5WIi2a+uPh1bWfp3jeJ3w7ljvbd0S3
JUjCVc6L1RlL5SAMUuZMXzt8Lg11KTkr5t0EPlAwaSfpWD/H+oiQ/wBaTiaL4CmH+94e6WrpsKgx
Av5oBm9UhjIYZqHD5h3AWUrnJRbtLHY2JYOFqIKg1rq4Xn0dXyhPJq+gMgUH7w0s+A+UGwTDI6W5
lf0A+zKf61acxlcV9jBxx6alslm4cxkONICr53JlfgeEly2Bz7mNpgs7YcQkLkmPhmGTKjeZV9TT
S9mkMnxl0Oc2MML7D/09xplIlm/+rptxH/FLPeT0SlxwX61NHvhFO9X5oT7CRGmtDOSQtiOZyuP0
YRf+sjCRpxC1S1uxKPKZLy98STkEp8J0uN6z6tiuOl1m60uAt+FCZm5WN0WqmwJq5nxYMhERlWtq
hZXske2KO/P0Zo8RQA86q+950RJ/fqZ47gn24gKFM0bS9jl0Su996B7tUCbV1SUkL9zSuB75cr8X
+hayUzKC7XhYNHcVWw4YD/vn6P7fU7gxIgUTLHdW9+Y3Y/VK31nlJMqFPwq0cUY33E6W/UvvEglt
QLCowqSmsW8vQtX7iqXHefdx//67zu/iL7bHz/rC0yJKWDJnBBrqWobtFG9bp1fRR7t+jGnU0mDt
wkWbygzUBuifREuGBbXGhGDsaG8zokVEIwB5cjxTrsshxNhHfrb38X8iEabFjCfiyyCZ7NHfAC+v
4elxoce59vGg56/fc3as/Blr5Kg9z1f1hH6Fl4wfaWyDSyRPd+Z0HKPpONVQGfWMydlUipr6CGPd
22+eUGfgQRG3CG/3EsqCjcTT8+t2F22yeqUj3Ocu+zI2jFFmmoyHHD9BtB2tX/U65pqu6QmQpmHl
cEdGpapWEN8Vg2xeMemW27iTZHnuKhHnbju2GmOXunnfpI5Lh8XJCexgJ82x7R3KQjCpBxiF5X+v
Fz3UR2OCi9zA1xd5/fGlS6H/sgiNNduYaDKa+hfc76kld6clk5M+Fyy2GrIuMl81IfXhZk/37CPa
1bVb+ScB4yeipVmGyo8Qr6pB60YwTxYJ72ZJsZNWXry2QVSCsQGo2qVXdSSgYuoMGTvYHkl0ScmY
A0IhGbY+Iahw2pEiXqVTtFT2Ub1JWi55cxOvb/ApMw0rJoU1a0leOEIfPxKmtQPMPNOE3s7CLzUM
+hNnHwXwhhn23hhiNjeoxq5Z9JdyCmhE8MT+h3lsYz14ISGdK5vQKsYXLlfHNhXIdZPzESjk9+By
NSO6897EIHoUBmIWhoSUaoJKcDbo/tiaQgjWpzZI+tphD6tL5UGg7t8VBpsDCCrpH/sVURcCRUM6
CpVmJ80Lk8MGDdo3RgFkMV1lT3vputIlXLQDNvVbJQ54YD9T4Eu323v0v2/beDCnWbrgtLgRaUHW
+NS1mNQRH0rf2QnFkmurIC+0NvCfc8Bn2RR2wMkcwZ4qebcIKFY342V2nHQHHGXtsYoj8p5z2pXr
aa6mTzAw/Av8YvDE92FDRWw0MrJzGdBNn48PO1pIdOp0Mu8GZkh8fguDcLUJDHtC3konOZNSfIoT
Au5IjwCONi7FNHshKy2dCOvfwImVutURFLjyA4lqL9X61LoCASSxc2G40Dd5y6/wm/3K3a+wrVcj
E/bDMAAaZrNx5nWqWvjIaaCI2xzkjAkxZ+2WsbBQQWwhobo/BKSO8cqQemDyAinlB0wOEjRExpYL
S/qouUql7AyX5YCvteDY0RU8vi6luZ3Y3sFqZ3K8kWOl0Y0KNFVeUh/vVjoLgKdwtQIYyXz+kNJ3
hR0kxrYQgfAq3ObOyAV9UvtWGWQCd2Xsow4gyqySRYZZ49JE6NVMpux3eMApnsDdA/g59Dw2GCJ0
ZqkIe+hU8xcfig1VEdRtIEtVl64SwBKRS1xo2+y1lEApNsFj+I9RkOYQ/lzVS+um5j5CfCjTk88c
uYepYzxd2iVaNAP+cfOvg9quLsECSw2pbVw+reLQbqvam+QQ1Ie6a7V3Wr2pO6PxucUzqLYACl0m
kzf+RqMZLdgTPuvXPzGq8u2Z1SkrJpvU4yeh9EWIFE9EulOE2Cl8hnzWdnuWHaQSuFqhW6VNbCja
LHPRrZo2O4EmNGi7nKXnxKes0AiwgZ/FCqYoWLwqm0+irIlyGb8DwA5m2q4jPJ36K/SNIGSVQgLj
ZZmDLh30uUzMK6aNS6RuZyYSdSYbHecbr1KXF2VXpj9wisgQdkslBqhAdGliIDL8MkUpt7r1zcUZ
STk+CmBBWylqA5fp0hY/ENbIKu3JF3ILnRXyUYU6jBxJXhSfeB76yRPn3RfMfrRtiofXdKq6/rZJ
uH3KPTuibL6SlewCgS/SwNr83SpEP58TPejFaBzsaPyH50SH37PcAos7hMMEgQZdBDe6ZzpCOrNE
3MECqPqt98U5Y+L8CBwRjO+/xvgnXodWBW2kajhxUghieQzW4vyq+eu0kegePh1v3kNP+TarJZ+P
5byZwMDzfnCo2mlDm94U+Xg41Ca1PJCQPdsgwUZ8fIkQYLJxL9Ryc0TzzvsiVp++3qd8xEF1wJo1
OX+qA0LXgyvP59k/HOjmsstncRs65DOJiMHcsptcomWAbSIBG4NWXRSozXGWpMgqrisgjSf7JQjD
noKXRrj87fpZbcFoN88p3j/4/TvnDo7YeIPm1OkekJCrY0cNpjcrfNJE3vevzHAC0TsmiUUiQJTx
QRr6W8zIcJ2DJpzvAI0XPKO2G+8ZxJoVxa8wTn472nXLVmEZZjdkrhxEJz1kA0oFd0pCXrhrU0Pk
HHdhCrRDEn9fdVrSarYNjaVzXFgocpUEs+j0HDKIJ+ZJghL4bCWDdGiffbQxlhWUhkhWjsy+tu9G
kP0PLdqw0P8R7c72Db2XgEag+ta+LNUHuiNDu+ZbSjmNNQypX1JPgGRej6A8WZWG5Qb2FxIdQENv
Up9tlgXCbs6T3PlgqTPhPmTf8XzkKln7368JdvICkoRf9iBMtNd1dBiP7TKo6LB1xCpFfpETKgJs
TKSJWaYb9HPMa3ZFLYLjWGYKiKnch8TS/8YIRefXNp+YDp20tpwtR6bo+vSkC7epsYw2X07B1lMW
p8en+p5EMgzvmw801hW45XzqfpYpR3AkFHqKeiJlYguyPjWKvzbl+4bEh2rksi02fVxf47bNmrRE
JDc8AEn9dql1cjHA7hdpQQJ6lHSqM2qGmxFl493zN5GNtx2zDCF6XBA4hyCaqgEhRD+wwXywKQbv
i99+u5zr7Zp3C43NosZpEJofNZfoD73Bnlz99H3QrM1DGY3Edakk0EwgMYF/U6FuruGqolc2k8G/
caauwXfDBNZH1cPIDKHDvYg4HmC+22gJn6fh5wAescK6/1TbE71KpDA9aY3/gbXlH19tulMXqnot
mm/fiZSNkAud6cFhWroHcwYz/ntIsugUpe73VxSq82sRMOkkLn4/hKso0iDEgH686ENT2SBxyiP6
VEnRh4ca4AUEIlUxFc7YMgCDgdNzf+jzLz4ZhczEvyiK1gJVAIk/gvRw9WZZxLKEfBDwEKg/zGdx
POnP0Aw/epMKCPCPOfiIF3LHXb9aGXol/a/93z5L6ltoGl6O7kB+YyexspIhwtNwqTV9XdrW83sR
ZPloeQ09Pu6doJvmTqTwjGHFKTjx58xd3h9hCfl3H4TMTh/x0unQFMTiluykXs+iVIuJ3Vrm3CIG
sSls/12wmJM4E5uOFJarrh/PjbonOz6xBhXW4AGYXs5ujnFBT05Ed5zr4T578dTyKoR6+/+IIeBd
ong8J2YeikR0X3bktaSOBG8Hs039CcOF7boazp8cAdjnOlMtp2SFwYMIZ8EsUHQR1K7ZAs/TcTVX
qCtQHwQ4FaainIGm6/8BkRaRjXjolqVZTjwFbU/BcGLD/igtM27k+F+rLuPs+/gd5Dq82rGgdeAg
UKXiglAMvM5bhW0lWaY+g8dtKiK/gDXRT73VWaDQUwnSJIp0a4PMbq6tffplsllikPTcnsLruXy0
/OrvFIl1tT2OXBDaXgRmB6aq48Ira/W3o8Md/Crf9DNgg/1+XzRvFsSz2wgvAN5/CCeFQ9HUgHqQ
dMTms3pt89ElykHfYLur65Ao/WTf9sdqiLrt/yBJEuIFabsZ2jWbx8pH95AGMoksVBMeg7iO1MQD
LSAC2fowVIWpAjIxebhtgBFB11K2oPbNqeDQB5k63lH8CskddDjZghV4TfClvRSTGQVaQTyIC+0G
MrpD7bQEggcQDdhE+F8OK700y7Oq7i20lu8Tok8ZXeZJWcLqZz5TfeNmbQmfjDIe43dUOqKwF94t
hN3sGZg48pBTVqVzywjcr01Ap2n3xj6RtYUOB6eymcQuTnXGguuGYM+OGj0XaoB6Qq+72ydiyVtS
7oWc5Y6poq+D9UNsQP68FxqajOdMKOCOmUvQjuw2IeLiGTIPsYVHGgxxfqsSJeWy4K00HNnsE+AV
SZwTLZ3eKIf0B7MFSW2dyg4Iq3hFbQfui61SGYCZTD0AN/8zITSGjsJwfFalAc03ISXyjBRtLTOW
r40q8kOic/fC/v31xi17fHE32UpZmfcBxGahNdwJvnb+8TAbqAH8fyA69n8C05Sggerr0eVOGSz8
GMcW3I0Mf2048GQJ1pgOLjdxF7T8Etakp9LzOuLc22es/epWgCfMli/8Oe/5R56a1gWvChfKz4m0
Heyi6niYwEqWETPHxTl4pVIDz8alkSq8taCl4szh9/dB1sADkqY0jFVY7/JFXUiKqkodttDz1iuP
3GqXGYE5uES9Ru46IWLdXYIo3q39S/pCmKXTbkkjtoQuejaBUClQ0fT/n+N1BoMs28As5EeQo7E+
RRVeylgctzrfLeoXSNcYP/33uC9IIBQf2IoHJ/reUQ6YTjF5gp7Qlbubg992C+KwCQQi+q4V9Bv8
eprIQndcEZsb9mEIkhz0eqO7EDsvM+HSDeW2PJ8trjLveg/5KjFfY0n8YhYg0BwVTS+As5g19Orl
1MC7gU5/Cv6I72O3DatL/bgYTRR/oAVsNVQMSgByovltuvHuKluB7mUlD6Bxz1HUtt21RZXpeLWX
eeQ8C3cGvDUWpk/CiW2kaVqrY5LPDy8PElMZg10vkuZv8rz0qCZumjluISjkNMqeNOFKV8Z0bVYt
WYaqwRbXhPTFm3e2/7SYJzMvbVuuivZ3M/mMMeI0BbYU+cr/Joh9l53FElhNPbtVy1LHwB8otFc9
vimmTXSV/DxMoA2If39PdLBVO6BwpOWzj9TG76LHG5VxWMiKwwU5An2Nys3NK8WMyvB779n0S2Iq
OAqm97+2tt5vCPpDbf+QxMBl6Qrw+iyFkKALhf2pbzdosDgxLQW/OVi0t8uZBUq7jpW2FWecvI8J
K+OUbG+PeI4+0932FUDhLz3Z20z54DG7TGKLFzYCuifchyT1Zd6oND+7bSUkpK9AlW+9b2Ro7OZ9
JYEPZa/lJfU4CLWzuL/NhPopNbJB+Dxdiwx3PUlXYT7Sz0n9Q2i//eWE/mbwFQErnKdp9nSpZhnf
o/CkxFhDCj4GFqOgnoenh31XJt4ljJjxfHMfBXN7v5eqLFcpUq+GNTqT+PSLdKy0XqCxOsVWC5n/
etzKGJxavIN4Sa0+JfNpcMEddIaJ6pEAXDup8BqYdYUC0UdBA3IYhMvfYJ/QeW8OHmF343mpW0k7
QZARlLGNVlRqVoH1smtIwrH8q04vnTzEsVajPOfUHzpI60yKJZUGzPBNH4vrpQ4vYzJJCODXWm/i
98h3V1F5wvPrJR1HpQ7FQUsb/BJ67owibkc9e1h2Krdt+bfQVnfJbjYZGnND/1Xl14OzcR8pmnLH
Lw2EWNH8LrX3s+/ffmUK6/PQp0yensFhM9Q1AYdxfyqZXiG82nSlcb7oWIhx+jgMd1xhQ5VAIxk+
kKOggaPuKbAbg0QczEPMRVtVYjMKdtlhlavxVDzW1iO9tA+pgMsUznnaJNQmN+aui7wcVwFsdr1d
K5mXZCRtaLRRroWPs32nof+Wg7L/X1RglHexpriFIMsawHhA1UiIDQHCRvLA+7j216AMSLf5PMDZ
MjoHZiehUCHsq9PPSmCpioJ2oDGNpBla+LBJSRHVReRCysfZe3b1CSCUkvdkw0GS3HCdJjAsKLMG
xquA77iOmWNebKcOMCxve3ZI2oF0FcqBDFqXHFhVWV9d968T5v4licA8BrhdrKVQzNQW2N5OPmT5
L+L+Y0Eh8nvfw0+xArcHnpXTG1ynvkjR3SGhP9TrK2pZkDtPMEgmqnxhLC2v1cwwRK8StNT8pE9l
0319ARSko4Wtd59FNH/TRc6D5q7iJMbjAU54EzFaraZDW9TFSqprO3EEsltdb7n68OThey2qRHMk
gNS3pP724Opdju+qrW/9/yzki2M7RifT1QhXtfpYr47usXTJazBy9N7KvTUU//FXDaHO5YX9FFLM
QQoNKSXxYlRUKis5Gz7K+HhGrqIheYXa983WRMk7paBib6Fc5oviWrHP6fkmbi/eXb1zpUmeXsCv
n68kNwhWgYddD5OLA3hsP+IF2CHVYtqXXdVtaqEB2p3sPjBpFZpY9bYmNtwQbx8Ej09RO3bJwhYZ
u0LZdngn4DTCDPzpvHNerugRQ6+TsjdzVk7L/CERhZGJVyuhInnnMNk7DgblMPBCeG81NXWFhJQN
gTt9FjpAOjJfPtkVUIXoFmvGQxJPaIwikPdnLJev2fsoVUree670AbI8eSaOqzVb1s03Pb7W+w+d
G2YNlJSCvz+lUkPhyE/SP1WzMs3Y1xLSJrbXLxJEd3LF4QN0+ZivtheOQUlONtz8SCEstrscCaWZ
uo1JaIApAHLpMcW7RNAKiS7rtg6TPzxqb16VL+MdF+8zK9MRY28A8wyFEc9k/fuWq4iY940I+uvy
VW41AxgTpE6pScGJ1qtxsYq2XiCLMB2QgwvoETs56GcxVjnHZ9M3WzHNZaLWHe9tODGHtwtgMfag
ftPhAIhuF9l6IphY/vxNUTVD4CkDqH5DQ8DajlG6jc90GKYps5CpUI6WwzduBMf6PmszHGUJuuQv
ziyMqJbyDuTZDkG3zTGaHTUwT0mMKQhW9R4CCTNPjSKDp4TGP9sFcdD6vptKWOp9Gjf1UI/2OC2C
Iq3Y6rEtKHO9iPBO1ly5l3zoeZ5djrZZrvzeBovlFk9rWRggw6+oogOsMa9I4JLytJn3dt2nY/9d
u08j+VvjtIKLyyAFJM8LyY1OwmNRwryY7GzgBK4inlEUFa8qk9D49LvnF+b5NfFDEtHbPu7BLCU+
Q2eqoPUVKc5RdPWdMwBVzOVQrAWMUo2lkS+i0Z20IcPGvs8eWp3i//CUeqOgQxUpojDpnwr3H9E7
BamUZtAIGwli+fxUGVMNM5zlATsurl8IpduxH1E9Wr+tgvPxQjgPyh+jVuLo3+1tDm4X0FHBZ21r
BSfCpGuX80pLYr9/UyizulQFe/I//ZLdz8kBryWX1IWBWmqPJzOIkjXe0AVjExLRZMnzVEy6ADyN
zOiPmTHefIiGqW2FaL7zDgNkYakAq4cqJXhpdVYkla6qjGt4mV/q/BddDri88K4+vN5JVVDsBviv
W8uluWuIrXm6gdhGTOmAoaFqGsxyIjadsQ0IIg6GCutP2QlgPsZn7EaVX+/Z0sWviPQC513sB09V
2QrOXWjIrka09dxBcbHHkmohU6RGx6sMsfMqMKTro+wBchW1ZVrcYvMtFd4WYfLjFdGlcjrn3Iep
QXnq2lKte+5dUVFA3JA2voXlw2CNtRMM/nFgSWIzbNElwEOkoMSTNQaVTS6ag9C17C/5eBTGISxf
Cx7vpK4imvJwBoZALHYlZhwJhhuXx3gjs8Xsu/MD1RBrowringYXeojDrMSLQh8y+AdNsE+33at4
cO+rs6XJD21fidy58b5SGkj7yQ9bD+NVsp5Ji7jZp5gI1Cm2ipcuUSanBIonI5bZctj8kGXYyVXc
8vwOk5Bf3/TVa3FWYV3g8tfWMbLGJE2bdg+iz7WMGcYmVjrCN3rh8fqMCfb1fEg3m6+l3WkIp/SS
a+GAhtaqQGL8e4AATsfYWzhaCV8GQ5t0LXLYxrD7x+uSTABnPyg21S/kO0j1r6bvslVhBt2rOcE3
wH/ShJtgSSYsIcSyL4pBaQ5Zcz8Pz5IweEmQhVZLHcoAX7XBd59LFbpE/cHbNvwnvvx/ezF+0StG
MsVMoKeBOKPrwccDB8sF5A8AE+UkxhrTM/i3TnZXbtFOEn1bsZIDNG6w9sh+7jP8sBgBIPBEtaM8
40DBkSLbxduv4ruGLWSal5EYRamuMmyIJssIY1M/TmqAFJnYG8QSkg+pzNyaTWJX9GMBF98GvCME
XRuX5QFw8l7Is+Oesk1tUWFpf0+f61DMt247WF5HoChFpwgiDbzxYnjH79KW8iv4I4f397wujZXM
PLN2spsN8piVpjL5oyimzD/IOQUkLbf+sW3/SRsqoWY0dT/TuN5THdkv1TBgY82x8atuhqFqxwI6
c6S1jgOdR/0uF4gtBSbz+rvaaH7+7sxHgq7DXwLEj/szDcvzKmc+O2LD91PfePwSJjR3gIN77aLI
9L892sH5POeZplzVdoPX7tEwH+JJ6MXQ8WtxXwCJeVy8U7tG2P2h9ppTrP/Qd8DDbRD7KzaWuYuJ
5tAxR0kZ4cI51iAfUnWKNEncYrecC+e3311SGTg/XfX2R32v8N07VJMMxSO6f6OD+DteLT2blpLW
6TteGWHlTC0gklSvnuwqp4gCtNGdUfRF3Vzi1X8eY4JDQToyp6F3GKEusa0rgOqcXRU50oB+Dor2
r81Z+g1RDiqQljG57fiGR7idUjqxTRYwOZup5lxU7yFFhU/0hAQTKw3SK5PN5gtYkRiw/66i6k8M
IhFT0n6OJyizWOuRvFNufSPiOBGAHEHJ/tIePtONr+sRsBwB4muCZOHNHAimtVGCP188qarBdrAN
0ZDH3nzH1EvD6l49/TCx9N1WnZ6FmKZd+hzo0yuIqBkzTgf0QcYxp04ZAVN3x29sYoEINAeZQILg
EcJItVXo7VhNElNYGJrclkBRWBT8B/FYZjeUyLCZQRPplnIXHty/RGZuE/vWfZeq1uSWPFeVfh5R
Sb3HVFyjobTU4CFrwqSnXipy0NMG8RF92wmg3pYN9HBuH37CvCoVPKe1p4ds8BpGsr6d9lTRYN6r
qM+8QAMeG+/TqsSFXnOQDYSNkiLd59fQru8yW3QMhHYdl6h+nqxaIk8pKjSJ5Tp9p+hHDbkMI6tg
aQYR9ZWDEYrtHLJDJicgiZTq0IDKfV2K5hzwWQ5aIalZOrRtLlSakVxrUDYGOXd15EODLQi8KvNR
Y4ZPdZmwPn93eRKDF3t34b9MdBxLmelGsUg4PUngB3SdQkmAX8KmTZ9GRDfAQToTouqZXpV/iu2e
E6CCTUQmlNKELzsVVD1vUfj0Vzp1r/0VM3225+dtCpCR9yF6tWbePnd21q79a88ss3ijrHq5f7Me
Ag4EKDUL1J9pviHbgXNaWHT0L26v6MF9GXe7/CDW9bQ6xkxRJSmCAo/NDqHvHbra0uJKV8u/NU8X
TzGcPvPJrIFHvRxsss7ATK/NOl7j9I7DjwpJwhPDDO/buXfEAxHFGBwkjISVwtayc22n2QfijLbZ
Z98xSY4jn4XCXBt8aYH+e1l3JqCBVmqXwiEvHHUpzDr0hKFSgqyTUtRv+NJ/9vxZQgTMiWRUMIsI
F079vjEFT9mzaYiSwEO6Sw+pkJ0avWorMA669fkMLMAb71dxaHGoIBFiRwO9ltcr5hC9OfN7m4Zq
xgNRxp7JPTWq2sdN3CfVjL3ogtjj/tzBwdowV44+6VyOQr+H0YT8/eubGOV3iNkyJsW2qifONZW6
e9LgwF0UnufUQwqO8hZzLfBA0mtaw6L3fBhT6hs2ohygCYA6S7DQIA7SRhNjhgppU1jUyxUJL00P
cyyuflHmXO5A93e5YOomz9ERZoJrRvabb2P4RGalo0TXUmkvGrDBSCFUKDS4O1jVJxzUAC0saC4h
q2HFEEQpxsoa8M9GCWqFTKcBryFJqqSg9Tz0kQV9AmbpgAh9xfipCkyFe4++BRdkVnytizUuV2vl
FeixrijipLKyZA6OmLDatgqQ7IfFEuCTCWWMYVd6V3j6jGQMKD+nMo7qQ/SpN9d8VlXwrFL+Z9Y8
x01rQu0pDrfCGdEKClYUBldszfS+e7FA+amoAIxNkIviedYlumtnN4Gn5QXss2cLUXUNawoHEI/T
lrQqZoj0S6JvCwuAHLKbVycDwiRjNHm4kOuAvYFYo0Uchbje2uI9EtDYK/YKPnDdC2MkLBvPTxdV
6lb8HlhLeECoN2fX5OvZPz/UYGPcZVfjZo9NKUQhANVDhrb2dRn+wg+0e7r0AenV9dSZIMCzdGCB
EVVm9WAnK1hwHFpYkBsgfBgCn7lXfePz/hqiHa4s4KP4/TT1bdGNYnJHX7dcLr3FArXHPRRKSqJp
NPwVjBLDflXi/c/lBCbwD0ATd9Y7MT8/QBk5a1ul8qWcMJMUGmIYg+MBFsjasiNZRlzJGrpb0B6T
Jnuy2CfzMnOx+xYIKUkldGuUc7ViceZ0qj2jX8CCDLu3WnbanVtR3gz6i5bgTvHPaYpUejZO9h+0
wilVLGGEbzLi1o0oeFSYNRHTLvVX3BLnQvVDxJYT+VymP9AJjMosmrB2qgswbOiF+bR9TBCTvdwn
FwC3DQAGo7Jnig9tKbUznxidbrGcS3zznuZidD9fPQMqe24jrEkowe7QH++PspZzKnT7Qh4mqNhv
/2Z6OJgBOPF85Gb2m4OVWGUdIitKblLnJvEOafLKz+f0ro8vNLv4pqcxgMfiZdRx93R2Ow1FdrMP
aLlpMCFxYIclA/7uO805i+5geYKs8qWzM0gpqky9z4fODwFPIhEE/8NQhgQR+0XndDhr5sIniIIO
OpfrwoF/HLZARtoHEd4tabFfJABUeDs18GM+rhnfECpaC7q3gvK21XpvdU2vXPAHVHu1jXpvUYJL
K7pEFRhrNsIvUjfAblawin3bZlFV1Tl164xkXwe+uvzNSdxQZrmCDDkPwPMg+eyAxNancrrYZ4CL
J1+lm9Ukk7eIIRnyuiy6JO+r4FXak49KF5Y4Gd05Nz5hR7vi+VvUWww9sHh0xuQl2mqUKGgYwb86
Y8Be1BhBnZq2qUeocGsYOSjYoJVo9sLYAckTdlWZDpQ+pqI7inLNFVLueeTAs4e4zvThNV2nR/zS
/56ZbfmEsQRSnKvfE9ibmaqgeHTp4wrglVjE02a0KR1w0b+dj2s7yCqKlp1/c4Lt79w4Uo2UO12g
oBNO6ul1AcZjGk//INE+ScXinzhGYcBHe78y+dic42GsIXQx8oKQySp9wgbQFL6PWu9+4HTD6L3j
TPz8w8ddeNjUOVpSJWquhv5AReqOKkD9WR5DC23alLyzkEXbdHCZ/E77wR3joU0w3+24s508yvLh
t7H4efI9/7S02I17TMT96CAVj1exfuyFhruTn5Xx9kibCYONBFg+SE+QhgLae2blZcXXnZYlYQtP
xhCLNukrEX0VdFF6YHgszvmFIi4pt1F1tOU2dnrklVsxidWx5mouRkxcfiA55X0fvWQCqhWO30RG
FtQwQajJXPsU0lTLKbjTBiCmQUZJMn+xU0TZXCwa1TFI6PzDRJZVZDs1PjjtyJ/5h0ODpxioP/ri
fpSnA97Z3VSFVweKgz0yrqVlPLem+WCLwatS1am7PQE8EF/mY+hnRL7nXzj2xKBwmFVs6YYkUMLX
smJppTgQtpPhzhGhP6/cJv8UbQ29lZbopTR7Jz+Zuebkk2GjsQzxz0LcGP4a0n3L+9D723o17rTw
I2WWZ5YK9FTSEvnLd+RBKqs5HGAlba3pCG33KUS7IfW14h5dn86yQi5kLedJvFpFX3rWeVdjQZQR
x0LFlrmDy0i1zMdj3QpKwYhmB8ulzUlpis5bQ9eVdFArrqEaOnMgZCaH/k4RKBk92g5EQAwvM6jV
jxEMV24yM/2Yd5ZEEvdmqvw7NgnlHS+cp7u7bsMuAzxQ33ZlrAl7zXrfpSUkd6SPs42mRIpC5V9p
z7emGuqv36W8ZvuE9p8AP1Chv1+SSbbrgmWEJzhUzXvzcjGtY6Tw/69vWYPypNOE22uBr18qd3gY
nzN4D/IJJGXRtBCeTD4Q+kjn0GHL9Gj5MeDVJarVZ7IOwdx1W0TiLZ1n7pBXgW8jBVPfi7oBLtbk
Khdy+1BpsU1trxuPZMDtZ/YBEQR9SVyM+fhjp93ECuXTn18qF7mVGem2zpUrs+jUl9AnOy1SMq74
+ERkTkLA0mrsXbni2tze3rE5xXGoL15SGEvt7JoLqe96NHNigsPC7xU8HfMezI1s7xGf/VepTm+5
7AGbS9DO5grzEWCZ8MAa+mco8c2kh7wFgRlBnaNM1g33LLUYyxDHdBeTLDSoMpFZMRnKRz+iMJEC
8jjfYjPzgtIFGwHVn2/V4RvYIdpdV7t/Wq8TwP2owWtk01SeX9CyP4e5QskXqm5jBnt6vaJ2mDgC
l/HzRPNaOkxp7MZIp6RBo+VCSeBY7ibFzUQPtBrlMh3hjJLt/z7kqZtJNBVZDQW4sgs2m0Zy6kT2
XuZcQuOOgwLvFzdKiL/+zxENpb3eQXZFjWQJLM27DurEKQKAu0f2Cxcj7TJ225qnPDgNxY9GIXGo
wTPiAXpCf9nMjZN+FwQUnTbGPiooQAh3swHhckh2D3iIlkK5VMMR6tto7p8+Z9o6hscX4e6/9i8r
IpESW8TEmX/upHiJM9vPKAOcpmYICf1V0/tXtgCKzgHOzGWZSCoCjjqbpDbgkJ56ibymZKTa1uut
gw7q/xWTTAZtqK8ODmXpFFf/xLJ2qSLFEpLlTmjRMcHLtTiTa+kaXTT9JTN146PbpcPfGqNNYvlZ
b8ICXGC8pRQEn4CT9fDQwutuGGCwJA0IKguj+fFqA8tl8si7XesYr0hMqjtgSDkJTlJW9XpmCVB1
KqHqbwr2oIn0FjOXPfnmuciVy7MqMTL52mKoKRtlaE8nezHjGFSbiLCZ7t/lLib5OeiaqRaCiiLT
9lpo9tgiXcEC5AKaX2x6Uc3mqKe2MogzD0gYnAvZrXqmlW92BY9b/IOvFUlvcNM+DYb1xxwEqx+Y
Wno4NMcg1lOqWGN2xhBxnjWUR47MWrf0+upfRRzcEAR+LDwUgHuPqQK0ItO4jMD7luzsPiuxs9y+
8k43dcyhqU/9ByE/US36WkVyfUyJjaJC6d8bJyQ8951D0HqDnZIaLcSB2Bdv7f07GcTx4/t+P4JD
W5uxm7ZkErQTnNMEznu/UdHps1LaP63Sgjgp7rJhPq4nCiTq++SWMH3fzxicJ9fZISeELeSwGYM6
yosyaargiEAl3w39IUiLCfVFKbZ87gBAmgT7gyxKUtdfDg7OYUWW5sQaAGik40otWjF2AaCiyKzf
itrpP6xGpqSzmgiiibxbhPCEuVFVePPUUCX/dxq2aMX4Cqe9elbMNDi1DjfUnecRFuSjf+ZOuJ/A
gQOteE+uANstLiSNqoSOCh90cuvdpgvuUq7h+6JfNx1DkrtdeuJZKi6vXncW4fHsBZA79cb2PV18
CrAzGpcI0/mZQdcDA1LF7YSFpv5ySTGzCyEcYj5arPD7q/oXy4+IhYjph1LrU6YZwMdi915Mz7Am
2fHPk7lDS9jHGdMJt+t7BXCL0bnlSV7L7XcclGI21Wiz+kOrhKa0LbMNx+dxd5X8If8yl4QsIx4V
Y00YEn+D0meGe16cgAvvS3rd56FcKxoUhE9mhwsFpp+Xm2Ld0heoAJW+5sXUmx1lS75dShHo5sSo
OVweunTrV5xqbFEWr2PYo4GgkokJbptcjOJsSkQ8NkoqwAsu+4E72z8kp6SYT4rDxZCc+BALC15E
WHBvlI38CUh5ahc0DBQetvi0OeTTeEpkYMAjJE3iibGZgrIYL/nHNOkSZJDul4cwvC3jEJAY8ULi
DvyshnewN/CvhIvaKqN87wtWHCSLXGY+bC2NwZYgXwJONXldi23XJ21ovEdHU7FUregBfle1/5vS
sBqe8GSOvN0ivu6IuwlsJIYDZpcAawN5y8kJB2/sRkk0t/2hkdbAGB/5phcV+u/KFmxXv8rO/Ov/
qUjt71f2BScSg9TJ2HF8Ta9GAW6/joFS3m2HA6q7+Kwl7BCN0wdUS1UNXY5GVhj9lrIg6IbpfJLi
UfIUgX3OB2lVsB/cOsxbk+8ulB351WyGtnOI+Vpdp4M6qEt6jz+1MpsnsEnMgxeJ4r+atSkm+1dZ
cX8/81QAqY9oZg9wjHfGOuHcSdS0FBbLm2dN+23/2WxR5iaz7f56Gludgi8cIvHeEKwNFjoI264f
hfgicVGV8/WuSmWO/4mWmgRDPtegqFG65/0rWORQQ8qYF+8FZ227VgxzeZLx46G5qFRrs2ffdJ1L
ubfgzzJB8Orm3dAUeyjGAmCvwRXPjuUjwp4P2BBa/AEeHbArlcdElsPNPCPmhfRtpOSGNt1UCkPr
dFr3+PqV04TA6bp2ThG3a59i+8aCYFBUjKJN/eOTQ2iuSysd1vbXybn6hDcc+KNKVHPjxiI5kh7F
6RwNO6HLwadltog5Yu6e3duqoiFqCWOpTgFsIYdgdzXoo9NXl3s+pEPdQoEZlPGP/y/q0DuqsuZ2
CDvhH4pc/QPYC0Wt+j5Cq0Yj7TKjKQc7JV5nGm+I9q1E9YbxmpoXYbpRPPlo9eZpADP546m/LUF4
vvtcOcUU9XcBAzNOqJ+XGDETw1y3Iu/QTlDGU/U6865mjksmsxfX/6kyfRE7YzKVKaOwXYazX6c/
qVw6dxR8gYm2UIglPluZ701yDxNxubTKG3WhoybVbrXJazYJ8slOeWwKdZOJv9zumIq45O10jllv
8k2SIKkCFMcjyowMt5o/n086BkQ+c3vizKVg7kdlaGXCfvtj/iIxxltIqtMDZdyyvPCTfiELtEmz
nkplcMO8b2QKA9rr9jMDsM2dvSFcYCRkRC0CYZNtunkZXuR+CMkPCHnMFB7M/2YTWid5Q5G4QZcJ
3Xw8bDoODKVgTRogok8wtCuUaqWovD5dCyQ1Bggv6UNnEmpMMs3SRlOgw3dTBBJdz4BYE59dkko8
8DGL25BMT6t6z9UC20hmxHX7SL7GQioVxHvkMjBUP8sSH/grYeWNdufkm8BYMqAnhLibELLcUCb8
x/dGkLaXUq5pOvO6dQk7x2gycdvaFBhbl9hirWuVWX6FjAJurhl5bQqj2oeeNYoOHqZKw2gUma6M
HanTZfruRvo+WXCEepLRHUjdnZMhyoksamlxT/aG7FcAcYTcj5dzhsJUNyCAXIXVQueCv26A4n2V
nmJGBALJ3zx1tK19CD83UfXtstfYGzFEjibh2f4ObFsny5XBdbJ+fl72/6RVg/pDObuMHYK0Zxea
RFyS+vsTVq9+j2Op0uV96bBLxrx/fOQZBogeSX9v8W7QQi3rHUMGKuHLIvloVZak2Zw2cj5JNOHo
wgRiSFinXqnR+88bSP0DJJtpmO41jQbhV1oroBVjDGO3upmYmdyBH5xIvmLVUv+bXGGHfPryUUf5
EvgDCWRwk1fRL/9YFEyj80lp9P2oRhqPoQXHZgXzaN/qXTC6c1LH2DpfLGujggdSV5T+i7tcRgrS
DSzAwYNN6XsVRQbKBOuACa7QLM5zdSWzYBLZ9MhDcK3sguoG0eLUsvHUTpNS+XJ34DdIlMDQVlr1
SIGOtQR0+fQBpgXJw9I0MwPXgFKTBrZS1enKq4qw0D39J8AKYhlnZUkSBZUKbBI+fV6cUUt05d33
UNhXGcPtymDSEyh+4q4e35N7cN20B4quploac97mR/DZa1JeD4FSuwRtCpuWj7jL+UUBgwKKRgxi
K+nJfKrEKZkJIAh1E7POzLpGd8qUdVqNewucID0LFoMGztdJ2jPX7HUWRWCn++QkzdIP+F0vOCLG
y6xx99z7ohtAqfPKUkr52m1UUaPVgWX5H7c/0byRV8JTQ+Jb/Se7+6ZbUZQXKDA6W8tj/OybmCw1
Cg8bMOrfVdq5CETK9nKjvDMf9uBNjJY6F/9bmvCMmXsyt+R2bx0tYPaI1MK+X42brO8mQRw0F9s4
bpdYoolY6nh2cqOiO9dLYKXi8Zt0yejwjbPAg1r3TtToEY8Sqk5Ydc0iLmU/NM6HikbHxTbTjXYE
PC9fB17T/loY0CuhE1sIxpyakZWKqS+n/lsUvyoTvuUxjjA4UTlSfc9yBRlNGZt6DgaAH3nI/q9P
CT6YSIvXa4pxTjtYVZ/5HKmRiWPs+WebLEzW9jFMP4KdcSl0E2tFWzmlLfyS6PqY8+d4OmiBn3YF
ItTndzpkRV4F4iDgotFl6afcAp8fL3pfhPgKztNKzWNHkz9RB9JvDwuQFhBC5fn659NJ06DFps7H
GyryNc+9iu0uuGBXvn5Zu/APVrabBGIJcDiKHFOh75EWoforxhJJsE/AShwuPuCsTJDF9i/JblP9
xG2AX6fXSnqtf92/KipZN9sIvQnX7C18NHM7zE0dlzGV40p5GL4UNSw/T9Dnlhye5mkTa144PYa6
zPD13r5jvYLO4tvqKrG4o9nHqLzsCQNWuEm1GMtxbIKCsp6uqkudzzZ1njBrT4cXLVXdNW+SCS/v
NJoVla/n/Z70UPAOGTmt9POsRWtMWGGVuKD08nU92JRiHVHnmXPq64mWoIEmGPsBRedDCDtyonOy
uh8kNVwFFW4awdADlMsGHd3LTE5T1fQSDAxwkv3AVrQzhTx4UlWdid7vXMWln9PcmxxbNC8dYF9h
Jcxst6nxA5+wORedvhQKiC/jAffc5G2CWnU5O+L+IRUWj6LyBv74Ljr92uogdaqBkNDeZkCqElhl
ldVJaL/GybVv1dXybGfc8kcdAMN+qoZJymNmdB3T7+G3u2gxp7/yhlx2HLHYIC7fAjDbg20dxLcC
gMU2Oh/QSiFczi+b3T830bbwT6hROcdWJliZKt6cl7pNsH5IIaC2TQ8fjziI+VbHUaeYvtIGnA9f
e0cMJh339geJGmPyWxZoTRs9lNttEUjP/pvkU385GdA+/Yh73x+KCeIy7WkHmKt3t8hYrglVBMev
i39rYRZUZTLI9zl7EdvmRDKL1wlZ7pAr8+abKgrzO7jw42WGSroaW3NMuEUZPoq5PNAPGJvJr5VY
vBq27RF/H7A+KJokDoeI8ZleSlb8ZNZz3K8TaQ/aVq+XjDcRTQSIkgfk089rrESJmLEo3/GX0u6W
/ecEQ+2sCA1akswEEEjRhb7Uzeu2B5eAbozH5Vrg1seHKDcCVsMx5Ull9qpM4lB0cYb+ayAn+QtJ
FnkN/ayLVtrY7pfhgqIMX1ZFt3KHtGg5t9ReWjlEW6OXSXGOgicp3BVcRlJ8axuzAduMiClsH5Go
6fU7H+OfQ5OAIBUwqzwq4XZBWIC5Kyy/WzO4ZsRVmpgOtIX90pwggieGtu13Va2RVwdIZLpDyhH7
49GCoHJXkguR9E8SHIRlV+8XORZCxcTx7YZLk87oLZKJZKrSC9GRm/EDiT9Lnm9G4+V0bpAWnCTz
Vr5EqNdcBnA5IDKKFt5oqldJAMhGRc3ntL938Y9O+/r2TcMzfKfUfDSs2JHI2uSrqgXKoPfmwfy1
djGScFZ9vPkMyhJvPP0tcMb3yR+NCMBi0grVIAgwKC+vg0pBsEapT3xXx9hi/doSXgJrMAjhFJAg
xgabIKcsWR5mDNdGM7ytHkAGs8jqhI7lIVR7xuzbp8xm8/ldWv/HmDclONVKAuLd+89DGep+c7Vn
Jxi4HKDgqbTxkz+hVNKZnQdaORo3Ugw/LTyW5sz6nGspVnJTPJSRM3utKbEFhSHGie1657fXHIeg
IzChsKAVEHnYsEwdbRskfmjFie4dEGPfnooxq9YRJnxgQmyTC+pdQ5VBJ3xDlkeQJS0MrltzajtB
QC2CsKzonyFy9UglZcHCVxIi88emLAU+mNeGqt7wKwd5+kzhVWwAZ8h8upvJUSjeSAGe0BY6avZ2
pLrCEInxNyov9wl6v+MCn5e/btIXzJo0Xb/D9/g+WQB7TyIYBz51CH7DkHF2VWxQHIVWgBuiBOWA
Xj4Fjli/MnmQWLskJ+S2YKKfUCKHR5q3HJA539Tt57WzYwmobIWA/iYFeAs/eB9npsco7pGMShpQ
9MBdO6WfEyW/LtRsfCpyh83ZZRxUWG+luJZRvPphbGl2YJIXkHPfpV9F2q4i/wqhKyvjtrkWkRSy
bS8gLsnZy4vasMAZcBz4axJrtydkmc+/+buvYpktuvuNTYJyAYVrB8Wbm0uFtUCXVqt5EUxKY/q6
34bFCDk8kyh4bYQX7VhIZWojrzvB0uzUFODxXysVg5pSISW33ocekqIC44HTQyxuQ/U5cLRTRv6W
w9cYrspWBM/RY02vuoHFkgZLzvOqVx3uITxYG5+9MQrNW4SPs1WsuLrKO/bbB6TK8496gVPAOAU5
53k9MrYlhBpmrhF38ib4dttebK6FJI371dOzRLjIOcVfdBfpwEXnHCMF6Cb+riCUQ7j5+tIKB1Fl
yRDpkDkHDlBDBYVvJT1I8tfhGiuZfKHJYrVSW5uyYJXPIjUg74B2Ka1GXO0mj6u74rKelYeAVMop
aNraYG8Ee1I16EMpRsie0sF1trk86b3LpuHNg3OGds8m1FzEB5kdyUiYSkcA7ZoySSNF33UkelMJ
UK2vn8X2pbMSCoIbpZHuXu7rrs91Sm1SDDrAlxy1MvWFiJA/hCea2gilYDAJWfr6DvFCYOGWyn6z
rR2CgD1NBED7AHq9Z/1b0nCD0VVje9I/Ecs37fGk8CaWWRo1J/eXURWco1SkM3+YPLFkM+178Bct
k8WTlPhzi8iDujsQ32xtihNdNwae5NiZlq81Kc1I7qVLM7RdAeehrP0aF/nvIF6sTxnpyAFe1HAQ
m3Zo5en59bx78SI817LIfoQ6TUZ3A7Cug++k8gTWSMlKuIf9HmVs6qIR72ILLbNpamKKZpmn+iOS
aXklXGtOyv3YAVDf6hDtc9a/advpil4LZnEPvSwcOheJI+22XPKz/ZKdwKaoaI4VqFoEK0tAYbCX
8I8g/ZzWR9X2yvWPMetYnp79E+uNIVzAM0YXn1vBaT9JOqpw6D94EuqtPyOVerY6EYfSGOdUfwmx
DpKPuXPyZM4INS0b7K4tWyO/odRT4PufpwHf6MiNBqu+quidoPLtHLECIGGUQkVm51OsrpVpPp69
oBXHjiwMenOgtJIKWgm/yZj4kkdWHTFC+0ZWg1CG2/9SNin8IXsNy9ZSSQ9VrvxZSL5rO3bM1sdw
DKi7JE56tjZKZdEcVYOqpsQfvgN9GPbn78RK+Bt4GMSQr86zGHS9mC3gHDwze5/j0KWHpjKQpBdQ
80amdvYXMz/3cgPQruablPYF2SJx9sOg8nKLNfO1kx+L0o2QVkf5lJCTTx/Xhk0PfuP6EqzQstCN
pdf8jix7mxH4KfGW9vG1nJpEzVsJNMvTKcUhsMWUb+U4lu58Nrmry61x3IDDuC3SADv4e/2OnSe8
iBPTky1WtMRrae8mTx86oQybBEBgY8IbAvefjWfcq92rv2aDkps3hF7SNPWU1ILUx0h8nlswj7sC
z8OiGY3GJQ2M7AmV1bRWwv/fxDaDeVAAj6KKFCh0kggbRcPeGxNHbUctrfXifEUeme0CzXy4jGfO
0F/EKtm4nEtlXqqXu1Qpzn5F6TAcf2q60R5EuA9BQGlk6ncsJcXGQwJTFH0LDykKOBDBGATxBTXo
slcTUGl4Yh6ywu1qWDkh7xnEOOXMqd9RNoFTsJicZOLhi5c/zplWOyZ/7CCOn8mGScA3j+2Fa0Yo
sIoXyccLjhRqVJavyNJ31CzO5YD/4yIJerdCgk1RdwAwl7J70HgDMVXMNY5wdINWEsayRGCDtudx
n9N6Txlc0wJ27rkOf8s94JdO2URj3tzvVkry3mTynVGd88zlSibHPrk6znN649y7/AADg6/3StU7
SoXxqeMyr2I2hnVwcoTl/9Yx8+NRZ07eVaarQ44lJ8eo8EaiGYdM+zzJV/gFR50vKcPQd0hXYKjQ
b69eXUyrNFUMPPRixkRFgVKU3pRfo3Rp+ENKSy+yMziH6FK31rt/8AZcuW6M8Qq124bWtLdqqw5L
vtd/BPvehVgSbfSuPzL590q0mcZWqXc1y/YNdZc3lRo5abT7Ym8vpP2cxVeEobUAUqDZNPSwoD8V
NQ2XxGfXR+54KrnlFTAv6hj2ti18KAxZ20TZ4Ux8GvdCn1NwAioIttMKG6W0bIepbccxJI6n96oz
9fJi6dxsknCDkBZhFD/A4Qbmdg22NSoF/fYybXxVOA2tVLmPqr7MnfxtDFi74GrdVQPLL5t51wXu
cJFu2/c+SNNL7/2ykgdheragUh69OAKONmAAEzx/O37tAnGbdITZWe03310R6blKR+8WlZeKxqqB
EMwTkXwjuJHnXCtlniFfWA4Dka4RrikRLAAqs9UMsodAAuaCVZpUybyOIGud5vOflsyZYjT+szrs
mHqtoM4BRZdSEl0CNiG86GrDMikBHcom/ErTEZ4NQUfQwNhPUX9Eye1qLCPHHAljIotYSMSdQXpE
MNEVAWVJzJvkeshrjMWSqz6YIeTajBxcHcR1rdr58Qiok1flM9j4VbcRG03Aapa7A8gQmIG6FsSB
dIweIhzkkKiP1eeQ5X0k79E2xnVDhWBEsL3ZKj5b7UOGkLExeUQy7KkUqfsr6h8qfGEP3g+Czfrd
p5oqSIbFFJjwe7zkHvPnIxLMj5bn9cfSxRsjSlCneXA4zz/fbLMwondmi87Cvhx2lTnK6wcvhfBt
gG9vzOsd1C/3wOI6FNRu0GXYnhrwWDRzaNHbjQZn3PuRuDtwMp3DNXODVcH396QMVI3B+a7d/+V6
1qHgF9e4ZOtr/qtdhWsCxzNOp6cDK0ObnIWcvXaST6u3FUQc4v1q60LFQJw7/Y6pnPqS/CYotBmn
oyWyGw4dY3ru/vCf84yYWa1PxOjTmU1vjyeug9C9Gv4Oy2UapLV5TghSVPCrD5vvNggxsvqnxpOy
xguY9yLmzc9dBsdjMJoYK1P87VSid6/MN6cpsbC0TIhHz8NwooPr4uCxZBErdSi12lu441p2L9kV
d8QPquu9VMZRjnTXb1qo9kHitL6I+9hOxO5/D0qA6JDhYFXv9IiO0edfENgcifPbyoorNFRkcaf0
JNlLLkIKBuxmfT0FE0FKHtvRlUpNkdSoGqlEaiKxmxdyoWI5pvJizNHfjtmsh0vvZaIC5HhqtJsc
HLb1/EMcqdnujKNVFuZMMNCmGwBoR2JWdpDG4r0rontj3AB2j9AkWV1LJJakjIY5wtVr+gSV8xjW
EcfsBJ+9ZvAIfOtkkK2oLFpYPnOZucULBFK/DVukeb3rqqTa7RKxU7+pZ5o9gbSj5HfnS83/YcLV
CSC/FQUXv4kDBN5MCtCPZAAX495ZkIFn3O7a00rdN5ieU3EmKO3ix2UZnbVKCQyzWZMAh47QiXf7
hOV3GRWlbF1tufaFpPxBkAFBsDK0Sxeq5Uu9cFfNEKU+R838f0j3BKqLp9CkKBNQgRhGZoJ21Vnh
M6sqe6JNPSwL3Z68aFX8MpjU3ke61ZVKLCw3YwpShX8YGiGpa3ctwTgU289VM1yTE7sTZxsS9pEf
XliHZK+zxibFbSpOehvwYC8ZofxBm6PcaFmM1NvrxzBTI3lsUybeMz8ra6fLPpH0oF8bvhditrj8
ZzMGTc33qYLjbYv8ZMEm9fl+B8sM8JnE7XORVfr0FHYHU7nGn4dd8P4A3xBnFvm7PzSc3wRD2kZi
4gdldc6CKWyPWUB6FgR8PUlH/j/TCP3MD0kq2tbDC6sLYflgTUAunaKFvrHTgKTk5O/7hViyi6gK
ObhmlveGL4cQTIA3e4z0NczgHz4ooxcyk6GA+eM72EjKuwJZGVnjs8nI/4dAW6VH9vOOIG5akzoy
6hf4Z+4T+6f3hO3YyQAozhk0tcQhnExJuSSSCSqyPtB9DCrXcXKLkHLNz7ErtVthzAyO+c5Y1e9H
bKTwncIkqx588JGS36FJdEYJrGnCwm0ypo4RGAKHMgRy9vwlkE8j5/H+RPsNCcywcWi3Rzb8cNZD
io+oKYJGVKHCsHHtrHg1C4kBeUiou4J3V0f5Q1yFzO/HSoLK35F2x8aaCbZXnwJfNrWn+mlL63E/
n4yHTzyJ7akG9NfQyol0Lkywqvpv7iiNFQm8IZXUY99jJhOvAnrhXlDqRVeHcf0RExkfF9dBHMjr
mYLQiFBl7rhv7lv1iMKjG4/GejnXifVn/hhF0RFix/gnC7mAdpZqfdl68Vn711S3T7IY2kucM+UQ
3vkrXctx87/+zLnHK7Yv3UCbKJPHdSHq94OFEwLSnTL+V1L1yEadumFhI8+vaWIuIbb8hBpoMUAY
llacJI6KHS5OrCdz/hAQe830+EP3pjTjpBwVwVE+CDYC70kbKrEnAV/Ac04KV0UEay70T5SDXKng
8fCrak1wiTwlHQfJjzT8IHoO7zq2IcsZ9O0l9ck2RP+NXAo+g+wmOzjzYit9s54snPSRwHT17ZD2
00CWGo5KUGxLIfKazVnh4GYz4v7VAiEvQE3BDzM6HvdW9BM8I6vkiFo8hzmz+tD9fHFucG0bKfxl
Cefq+rRSouMXt4akFCv48W1OfhKH8FvI20BkPo5+Qc4Y9MSMBdKc2/rDMatrPJsPrFbQestcT1U7
W+l5kYC/l26Y9Mgx4p3r573iDxPK2yYE9x9MfZRgdPFwF1xrX6tfT8q9qWCXSS8o9NH284RkquIF
v/FmWjaIlpciXbiZypDEw2Bc+CszJnMS0//iuLQrUOTZAH0kI/1JkzlMaZ6eh97NFXpp5pimt4qL
B5HW+uXzijV25KPxnUqPXlO7IZ0ZZqn2zeOUB+sphO9G/SHXyTttFRTEOswKevttRKbEJRz6ir8O
5QNffOGOVyv5cTJeYN/6UMhvy4RX7GEKp8e0bMIrKFfjxD27+EaU3fxRBlNX/4sHSbJKfJTHlwgV
XL5SRaDEXEA5v3Ne5BYhHiHoGIiYpa9Vb+0voWCLTUKoFr1u1Yxs1RC+C566BjKkuC812ShXnLkl
/1tVZ9YOrnr9lXZwCD5bDjALy5cw1rLXxPcNQ7XQZDY8GqgIUTXcj50VVu6+n9Z0eqCq4dEdoVrO
2ZaazH/SyVFfSoBUFskzdvt5o4gn9eWLOBZYxGiM+tvv1N8jpB52Gzd7vom4oi+Th84CylbXWO7Y
zzFimUlnpMp2wfbuH0/wPOEDqWHJBcIoDI9qx8gXj7Y3tms3Yk09PdObObnk70pQ9B8F/JeZmYFF
m/MUwRr5iAcHL+RCguK+r4r8QhcatWrQ+Pf+KOy3hFky4pXd7UfKMCy8U1HH7P5U3ZJ/eNDlP7UP
Edygh18wYprzSIoFSeWT3T5ML7jDDOSZEcB36BZ51S5eJaOcCZ5QgSu8kC6ldBuEp/C75cSuL/1S
mCGBXFatid08QdbOVj/ajjjRNQbtWj0fpYv6BSPgwK/tvN/nbe7WVvkYWscBMo6FMxCP0fDy5ccH
wVvlpLPbSiQTDxTJ2bKmUhPvicCsYiYwOD6Lxc77QuP6cbr1EAamWooYeXcYy/s/K6arQZeDDbnR
y6j0IFHdK4e1ZhFySxjGPrznfgBNxxjDg4mlnVlL2EC4dnVKoKbMWMDZFdbV4Q5nD265ZNcB3qLO
TwQnt7Nm6kybwfOr/avQLpj5JTftARvlMYP2zPSa5a/NXpFzOz676h289hB93ME0+E75aYics3kT
sb4XKNBmguGjO2X541vsoiu3M2Tj5OrUlDiDuS+TLS5/mZa2K05i3g6zYSm87JE4KMoOWW67HR+/
cYgNdMlbFoy0O8V0AFJwaN6BFooPhHblBIxRQL1DBAsWhyyhxRuGYFh5Wz/Cjo/1bfe+ZK5LCXJx
ACIPA+HJxICACcECbwFLXKmUSg77n2LgciqNuSLDjv/JIPzAXBumcFgE1Ro47s+GTwzo0BgoTd93
2s4t2xGVFHG7q8A9CAAAmlyy58HcxEwWAVQGDuXK/GgU1K1QctHo+ZLhN5IowVN9afo4ZBgzlOY8
pKGkKwbJ1izW4y88cr9gH6IqjE0VMa0Iz4Ai4iC70fg2R72H+9X+grkPSsR5IOvbLxqvU/t7RZlO
a6b1PfkV3sU4//nSo4rpVqc2oeNLu+X1fSyUTC6wmWau0t/MBTz+SIlypfLSDn/0RV3QrjzNCEpQ
j2qdXxENjx9vVl1aBPGFg/o2R9qf4G89sjqvNYvC2aXIo4ZkVhK7yfO1d+P1kIkPhfRZ9IdDYkHk
f/HqBcf+fFXCyc0o8Wn+4mXxuDiCmLfSM7f6PBNz/pKaDKvzIiB1FRVF0yQJ32pk0UpOKWP1NpEj
1SeI7tIpn/o0/Mwc1aoUR7bsCxZPhKuY98cRNTz56oU4H9lTZoVOYsRdGG+3Aeysla3f8zSWtKqK
tabyEQ/meCP5NzxGdixleK0vDKySUstgnYPZKNxHX42qC73xxAmsXcOXI2f+kuCxxSh3wXr3eFe6
CTdriTyGWW9n7YXiT0ogPJf0oX7uxF9HpUuQuODKXDQpwE94QHjD+R/ZuZSllaoErTC02RxJMar4
y5gsnfFPJp6RlzLUMZqhdprcoNnjbGYS6G6HnhfIKGXBT91qz06tpDxVDMWJtHT1UtGN2JkPsu74
8tVJKaWFAZJcR3HHcAloMX6V5aj+ZLL/yV+j43ZB0mDYRsQNgd5l1TOugnof526L2Gb+uGBVyawd
g0PZXpVL9D1lNHaKoimUtG7aoUXSFcscc2JJ/70/36AvcrQug/BE+sl6IMGjR9gdoBY0lngTBJ0J
ZdmeBXq9zc+JJiwh+1tFJ6BXBdeWN9Pw8kFM0V/CuXvVPvS8t1wH50xFMGjadwaq9n2UE1YAkHVG
02U5yAsUBkmerVdXHfG2E6SpjMtMKkuASUcm/2rAEb0L52dKZHnK1wmRrDhIPqxhaCx3TdhF5QbW
gGTMvGXwOVFhFB939aHLMd/NQgTSW8MpEwi3leo9XVXmLndyzhjeHd4sOnDtfvaPnPp1Ltu12X9K
7mGHnR+5KxF7N+DmkNxCurTaOuW6fayZrDbxrpMdb/IjiZOSmHWHY8gsrxAUc7bDM0YQNkDiU44Y
+M8K89SjPpbSSYaBxZsKgB14RCEPTiphjtbvGv6AOftJCdGNUNbLYEXaTmQUiy57UqujDh1geK8c
WS/rFFZMla9bF/nOKKAWUlTrF3sPlEl6gft/gXwxqpuq9igcC/+PY8vpesPim3LSEC4I9luzGAu7
7SIOK/dTdvzZ2aUjehYVaWd/7XRbC1PYvrLxankAQc0LcolH3m+yNJdyf0Clx6r5/y2UNZwvzn5T
12iFCseQYbXwTsyEKv619ZR0L8dOlKFDVl2lm0XLlZcdzGfEiZNtLyWx9/ibwcHrr9JSO+qkkVuV
+e7rar4uvCNlu8ZSDTutKkFU1BEmf/Io1umwO0N+2kG7aAEPDIAdPOsR8yDTfne5EdeYMdm/7nwt
la7oytG42JeIj1bivvchGH44ieGOhquixWuziPzltanEc3lQcWrCPc2NuACFTBgO7g7fFIlHNacB
DFyMVwk0Y/jJ7XeLmSH1QQvaUT7wc23ym/CsJtFfiEjincYSG6ZBGTncbzOdn9YKfs8qKeIFnci2
AfaDPsEsdmvC/sFFNdiZtdeA7CMUBf61TuuyIgo/OnKIRR9aW6KRXtvx5Uog4Ic1PXsSbNSJbUas
PVR1PTv3DGh7qfxcrjMdkWETj/po7y89NunOv3KLD9JG/IRPntNLXMf1HXG9P5Xuj95IW0zTDCMR
x1RUWiQlp3FkpjhEMau8ffIT0WV2PpQ6YZvNm1IB6vsM1xNsddGAxyxnGxLghPeS8iOfp88+MrKS
trBqokkR5MsmevEFnYxy270XqmopmGUk8nD4YmChnlBJiMDrcMHwEYOtEtxPr2JCkpHscZLJFupC
DfGCUg4My+msHCrGszMe48VpR0CQuEFdrBWDKSG9BEFkxvm77CVUu8fXp/yeuoEHYFfAJWsrYWnZ
Vn5Du0nQ1tumFVjj2UbV3tFyHR1otDrQPJXamTA+aTGtihTheopu9IQZzw/qGuykIZ5LiY1wSDdE
eEP87vDRRufjzfsfDXXX3kp3c5pncTXa+RPhBqBXaygYNGTu/15qEP21aRMItiBBoBOnZsVBdB/8
aotxy/hqvZfvZNxS9XoEF1bhzalIUWtSdPEKUhkEuwb3uzp7IPyWTYde46rtK7pkl8wg3hG0otf7
jhzmqOMETZThtYo2Ztz7kVapMWRYcQCY/amro/YJWgMuq66D1IJ6a72iRaKbzGWeL8nOL3xoOneN
Gi+SCTXRJ4RaGph4hlqwSjN3PjYZeKuGeY0rc7dX4NFnnd5H9kP1GHlb9eAXY6eOFvaXjGzYcU7w
tso0lZ8gyvGMZgUOesyo+DGa5+W8mdpcg3YklVKKmpHCNuYUgedq23Zc5HMN/Yxpodl+LD3f6hZH
413YvNoxPQGtC16U3+ygLWpmpXfwd5Mb3oMQv0GMNbzqUTp5BSoGkM3kI6TLcOQg0aL+E6DxR8Nu
mi7qcPJ60e02U/bqCwMGj6Q1B+LzmW9Hir/UPj/187Txljf9J6UfD3XJpU/oR/Irb0gqep9hbgpq
pc8qj2nlsjjTSbhHqd7iRNHuAa583M9gJDn1UvWPWraPy6oqc8KjGwH5hI5CsJd9uvhwzZVja/Py
fEI62+6at2BLDiRu86bm86QVh94oi+VnID/ejgfsxEkOXeKFrJ48CBh68FmtTG+LkF3VJAhe5D0o
Dov44yKr7FW3z/FtIHZ69oXTj1EZS0pSOHR6lagLQ1PWe8GD/5nY2NiyeLBbYZvmgCCk5YVXTWLr
GGzqG8d/0hmQY1bQDPGlG2wX+MnVpbgZy4OtYwyK6fYIPWOTXGJZnNDdQdQWSp1L59w0zrYvA6HO
5QtQkWRQubmFZkOrs6V2qzW0v4tpJ7Q4kQJcs8/djjdAgbHFCM0F4U98vrNSie2xmkR3s3tCu4tF
4jwgoVewFXlPWwioRPoJ1szSPaOd+3mX1GJcMw/p6x3OsUGb6o/0lKHh3xhDKvAb81vcTCtBaOU8
tdXBlWdhTy63MOvE+QU+CQUnUPD6nM0AO2BZKCMv+en6nyf6hY9zWq1gENL5t07mwi0yalTbHOfj
5GRzHAMXk3pTwHIr3nPD7QkULyW8yFTCBqUmkv2VkHFZ/2kUBjGEqivYoMSMnfwGNKYNXnlyoL8a
OCuGa0SmESASBeE4FJ5WwcTa6LcP/OLOBBPgGUu37fD0mck3ruPYE+Rl0doAyqoWPzezSXTE+Apy
3DUOYskP697AXGFQzso30mxRH1C1dQcKbS798LbY0cOWMqlb1tGAOL223FJNnGDEk/hpalRzQKj7
CiHQusn8F2SWjoT7/xuY9cxiyNA74SzlZhn2Ehh8VtbjNUD3YKgZ/MJX7f574yLCK48tRqfNsRR1
QXf9gEk9iwTBwjieMXdvJyAcvodiv2TDP4+6GAlueI1AfeXDfKvNw9s1DZ/XyqoZOUKfPydZ28+P
Timc6A0PKmBTpmM5Md+q7gKArgXVJon10aHkX+Uy6WTC6Wmy5BCqWUtvY9hT3lgES+zLSl0B3xDn
8/RH7aj1+kJl6W/1ygvxgub6vv82JiLHZ5A811PFnhyxZnVaT5+i7QIRm23/5tbBQ1J3ZQxpdC06
t0XexI7NOA9yUa1mHDo9ce7zcm2qn3i9NCTHqWA3ySw9eEFQMgROv2sI0dffFQmtVyhyKBAQhQNF
qkibFKJJOB+OEp8jAS/uS1xNW8N6iTel7Kr/4wHvAzyoKtEH9uLEQ/zHWNrt9pnV46WggolwFwMP
xxqdFbVwB1lOGIbTthRSzej1lnEX1iz08lHThG39LnZd8Q3loeipzPIBzC07upZpoFe4JzuSfkiI
kuTNG1Qd2st4eKM2YtioKjMqWGoNHqtWQObvYFLxN7SQA5PFay4IyhBPLz6t7D2Msi9Q2RhY0oTH
nwinRjNksPiDc/AovKsckvR8kDeXS6esxlRNeJFSY2rvmRZ3OoJxoYTvS/SQ5tAYxG/PCf8xdro1
KpkmgkoPbGyRa7FbMJdWxhu5cKBV1YQc60h62Q75xsb/yfXRd+Cqm5oMFcE3wxXgLVwGdzJ9S91s
/eKyzvCWp4M2XqbwYcs1uWzLv194v1LVomYCyKrlG/r1CvNkEtfqTeJQILxw0nkBW7tAHuvW4ZMC
AvEv7C2AuZOs1MN9BHTdfdj8DoY344xvYStkma1VqzSykJUMvLxR2Mnq6wPI5WhnkLRzSUjjqSbc
6dFhW3+t+4XdcvMRXiDcJIwfRmz5QQaa9Wqwt8QDGM6GEbl84Aae9Ke92W78EBBq+3U5AaDdF83O
OeeDk0Sb4Ta5quH9FbpMNTXzyrLBonYsfLqCV2YDT32Frx7il7RsUZURhJZC0kl6BxZioxoiUkxJ
HEQicB1PPB1/NpdrUW0X9LZdZdMXw1jq0yLfkZFYDmVSNovMvySzOnMG0uckcLslq/S6sbiNG38g
NExKvuqakF6w27ZPeicYx0RzXm3D/EFj5NEIV7Uf8MY44+8598Uy0hz/DMH7AfujVCDTL/kljE2w
WyvdOMiId33At1bDVz+UEOLY+tWQn9UC0x9+PPis5UQRHtXFDyhTHN2mjwL7ZjZ2/VO0ogU0vfXh
gZd62JF1bkVBmRoMVjkLH8gL0EV6ycZdmsun2fxYCu3VWkiAlSuyWIRT2ykUJRuMKg8lmD3oV1wE
cgZ98qk9JBN8V3QJsbVrq77tXEqRsNtiVAX9TLnibZQ2r3LfgX7r/O2ZmQtHEHxnpIzn6Rlxd6wg
AT5PoSpgDV70N98+yYgyd3669r+Uz0w/kWSsCafeRS6WAKr2uHaEESJ2w+WtfuZnQSxa3xDAhInS
nwHLIziIrDBF8qkZ/QFnnmX3VVYMnvz8M4/t4weZHnbLfdp8+QaRhTdhO69Q8u7tkUc9IxCoMGaY
fwvn86r83bhe1LrAdmmmix6dc9Veg/aO4Ikd9Nl9d1wG1y0/Fstzoz6eUvoruCmTG06bqsUUWMLJ
QcGc3UVBKUJv64mqla+4HHlKUVQ7W02KD+9lfaf/cONDVM1W+wKuivWqUNybBkPh09CKFxlDg6tK
7TQH+zblk0exALXSgQC6ULfNFniVhi35eG/o086sGOC1suL5s/x0kGj+IsjkOZ7PwoSeCRdT/HTS
Z4cSsDa79Pl/EmhPkS9OTjkUWMIrbyrKTbLG9guV0ip1rp9FvJkT+TS+3sfQfsLkgM/yqrOEuVTb
5O0NhJOAMU40pviZYBI6p4MHDOBfJa+nXZcoUafJ7Frgnn6PxNgkI/9o656Yxe8f4HTUUQvlMxYc
eKGut94EGlXjUeWOu5hRWgmV1TR1KIJpgYU+lIIZbtxswgf/xBLt0PR+Vyan//COkSpQHRODIMfr
YubGvYx2uO2b8Td7OiC2/D4KEVdEM6KWEBCGviToWNhIxW6YzS6cMC1S7BEKrWhyeYSXTQqzeUhg
B24q5MSBVz4WEfdBF89rfS3MFP5EY4ddm1xCamm5fjWSsf2DP4ogBX6U1n53YXqSWJZkW3TG1dGR
yC+oY9dPa5SMNvC5rQYLmsZ4AhwBGWJ7UbbhELykS6mHc9jfaKVIuBGW3aIf6KI+p9lg9oPGsLQY
0Alc0LjbF/vjxQdQONPzyLx8EQX/DK1kKGs2hfobVUvUcQ/OFWirFvE1vSwx2DuVFX5YVGTfYjIR
KhqO16QtoiP1eiVGO0oqb3S4lyV/V7+GE13P7XL6vo4jewVCx6b87ZiY+U0is2goddTTp0Se3UQo
c0Vsv9n37VdK4t48YAnvoUzUHvNHV2Ui878BkStQcgyLA6Q1u2Ma/z/PlO6taJAgghbGt7aql/8m
tFbrJmHtMon8GcyJoQFFAJvcHo9fUgRAJE/tMSSOX+pTlLGfvkNBMJylcETf9wX/MvpoTPgU2KDg
i4TOFl68u3ORuCHAhJmy/0L+PRElwfROdSMn3ABvJM/P/Kg3ENpLHaHCIrBein6K4rOAdxBMAxUP
reaAhNKhu9jMgmSpQBpssIdcUNTFq4PSn0ZDdJSrU/mpnJ7fU5KB9Qw9eaoVIxT+XXOFzFn3T02V
XypIjfFXhrWYE9YVl7c09GE4JCOSLfq2ceNssn519n7d/OU/tQHbSSQKTRUsGb83Ndc+tMB+rkrR
ZNOsOhMbfTU4tIAInMQH/mJ18qIHpdAJwu0B7G01CnyJ17uqr8xi0ISoDWqIjW3FaTlxLpm/9/7c
YOTGcYFZzzedpmSYh2LLlN7OfoXDHVKSgRYE2X4AxpKjDH3nIL5o8nNH6IkcMrG8aIcWbjndVUE4
7AW23OZzu1xzhuEGvuBjbX5B537FSNJuyGTvl+phjxJAOtpDtpaR8QR+b7wUNJixIRRdg5cms1JZ
iepoC79pGOQZfGUfH37wno2i/sW+vkI1RWS6ZN18AvHrBwbYekH0X6HXDvJg/ByLI7n4/yJwbtRf
aDWPtlt8vyB4L/qDJiAzxqJOWV5U+1WnA5IA91j5zMqrjagP6jax47c9PeZa51cPV/3tNvRwVHrH
/aksfMo65B6TrTIOaCRWM4T3K+JsIOVN/sAX06LgBELSfnJbOAEJ121NyVo5ujPh7PSaqBebj12k
/XWRw9Bzm+AxiosQjkWqucFmzqbk+n3cP6f4d7Di3JR1zVL+DWJ7luK6ApiLwSyWwlf729W2Ybqq
Z5VL2C+1lnItm1Zh3UfLitZj69TSBhqmV/+qLSu9AgvRV3U3lIP/0L/F7Z+KTeNBXFXN2SsWeXaB
QfNEzQHHMJehym3ezD9XwI7VfsflMSnSC6cWFquQYJxwhCJX9Kbek+IsSDrVuSal4Z4/Y7O+UhLD
sOmpR4TKLI8ocS9NNUT9rOMRgwRUCJNSHArn9y08I7yhWFPZtaQMOCzksa/fkSbPd4qh/KTpeqK2
fEDH9YlHzesl9hopL+u5ktgr4uJkajVbTfLbAf1Wu+WCyV4/ZrHAPXGwEUTcN3k2StcwgioVDZLH
TndZP+gQ4MbHYKKzY0ck2q1G+tKpGytdx/Ow02lgUDGuWW8QO1Kc24I4UoL2xIlxaqeXzpM+C/ne
eSFrnHY2BSyq6tmnAjkBSJaYb83oMkZQ4PTvY9/ubY2RzWWQy+8GmbShYhgMttYxMsoOOqvTtd0h
onghG3pN/YoJgLZiArt5gbkNDyNJCS/xU1lm2MGr+Tq4DIM+fdxvNcDqje0pYm16IItWIOAepMJl
OWOGw90TJcQxjqIzbFN+EchlZi6IJcu93xAhFPSBFPb7gw7TUxTIPBjCQ7Q1Rlv0ZyUIYtqE7p76
s3t0tBn7+eDS6qnHNFS+p+bCqAN5SqILgvuYyxtfE8SqMGiF8bRgBpHIsl/KH2hpNNXqyp4+hj8O
pate//Z6YnknOfNSR2TSmE17TJ6UOomAgRuwS7ycmDCZx2g8HlHmzoplgaeAJer2iJq8bK1K/lED
VrvcR81kCGWx55HZnle1PZDUXlgoWimsu/xrzYrVjQWIQlgzzv8EHXtJgqPGB76etAWybJEFXR78
8n40cifMWC6JbewelBBdJobaJlYhd28VaE8H0qkbe5c0UAkzbLoDk8SapqwmB1d4kL9JYQ1u6NWJ
1po9pDHOsckkNoTPOVQeKYBqVWZ6NiXuYE0MxywdOIh4jdbGxzKokw5fqvYKY+f1XUw39sCWtyVx
RivwIKId4E2dLxiHsmXlCa5G9KM0zHgNBUlqfpZqjK/WJqXQ3XutEtmRXSeR5FF05bTXLMhAATpE
n5PJTMkTqa1X5AM6R6MbFsxI/ATwc9cPKeAtG2pIYf1n+M8OXVI1zbBBlBI1VN30MS6/7+DukSLv
48YElo/fgwz4VwyU0wcUWBwvuDRoSu68owwNVOfD9YEx+2M/DwNNIrDOjDIUAgm9g+jtoCDeTT92
a4m4emSMxgVju7Y+lRre86luHSoRY2NPQgBbzV9pMhs/TeurzBX0j+GpDnwAy2ObtfbSPgW1QKpj
2pUdqvetxsXCAItZQQ88hIqXmV/237/BKzQDnitSVVnYpw5jK8HSRXEzc/kCkZfBIhfxGhwL5OLw
fYfiLdjRGx4fTcpPgOcxRXJehqh9C8PsHu2KoAtv8emOAyYsCLV0me+TL+G/G7y5P0A192H/0qDe
TLsBCcLqxdbCF97fQRJmIc4TSeRaeah2urcmu4ZRfdEB1wu5L+RtzKzCNWfxO+6jWWBcRBbnn79D
rgjMyoJVsgm2m5OMaXCOEeoWEzO1ubxtgG9nD7CikEZVjxyXNfH0IqKCTowBehTz3t6n0kppEs9J
IAy3ebmig/dSRYn8UndeH3CQexGhPy4njXpVAj3nvL6t+cKob9LGH8GCnOQAIA/G+QEnBCP39jJM
IKjDCwKaU4WIQ9E2fWrCw7m1yckZE+778bkIkpuCpXleLkk88Zapb8SjDXmjj/qNxcwAkjzdixKW
hD5+y9wjtmpre6xsN8LIMdC/pM1eawGghZ+ckBF5opIuEGkrr+dAGPW4dQ4qfqHLsPP2wLvvyOJf
6On/nLaPBuOqD8i13nCXWPUkoiUbBbRMAqfJINtUd/z1BlAmYkPLsf5T42JvXtmt07xamU2hEa+P
GlgovcBpd/pVl3d0CBC3S5I1dEz/M6WeOX667/Pb39Ot5MuLtL++CbbQESoIfkX0CPl39suUnr78
eIt+C1TqUbFmefNK+a5RaTKGPgW2wHqDb9pSZU0nfrllAenRpCRb7BZjc090IarJF89T3WH/AHAL
uA2pdpzTrFamnqy7kZGDbk8mYlzH753SkUQzq1WK6Bl0sWm915vUDsIoTOB9uaQDfr9fbnGhZVI9
QIm7RvSVo0hcfxiVt5Ww2VloVnnysuCl/G/e2Wtqixp6evrRUDOHl/PVBUdGQdl/MpJReOSPtilo
X/4Pbfe5W7GCLzT2dHp4Br0a+mHIVBVz5togJi7hkyvM/IMGFIoTGOjRUjD9MPH4e0pJk+yQLudJ
L+deeLOjRmOF0l0MT6n+fXXGKrEFj/I8mnp9xE8uBZObQzEfcGK+FX8d6pCat5kgStZmlm2okc0R
o00ZX+eyv2ncGaQNP6BVKapKMoxOfOY0UTSnNY1ird13LmykEw882Gw/e+44ypAD6p0PrsMehxrA
H/Yy/I1AlVWNjAfQjlFqvdQg1Ri/7UuUBYaYxtCCaYOAikh0/uqq+zPFzp3+/lQtAnTx3X3OWwwE
Tc+/d6ag1FNz8IDHYZxAeK7lhp3C7HmHK/cxXMeIPIKi15kZ6g+xlmiMuhlm58sHGG8KvETLTsth
OXUHfWOThr0kroivkCKpJ9fqIuHXu1eDlbedZxupN/7b885i2D9dTA3v4zSv1lccH2tGpHZvEjcj
LMEgL/+lFCJVsUkhwL5gG1KEAQdHNIZJuIDd18vSmQoQm6GPE67ZcZvgZAjM03GZEgwOlTgW1oQ9
m+2KPtv4DAowW4sG7gqKKvJ9riqctPBYaU1Ul4tOJCXQSJQTwYfAErykHil9dG7uWFxwOXGi2a2r
8r35uRbX3Xh/EiliHEcev7DzVfy/tRrfbnXwdFP8oplMlRCgGrVWY9ool/Bn6COCcdMmPxLEx3MG
LaE31wUVK1N+EWPNN6Nr1YqjLMqzwmn8fjJOCgIHUAHn+o+SDz9fxe9lVdasJykpYQOmVSXxeVZz
rvdjK6N0VimP/HcMxvIneWrUwyQDO60d8F6GQKk6r+p9gDBGMSeBNmdS7aS/22/hJ1EYsdNqwYZ4
7L+ag3WxYGhFVgtKkBzoGxXfA5RBpSFaEIv0QuhB8jVIecYNbeHf0P0oOyDVx7ueyrQgKxQyTM6x
lsZgpJMqY1Koqe88BhVXLQCsMdwx/G7Gbd2jnk0qPXHnXx19ri3fRY6YwGQB1BHeEBTQnTAgG6oO
qlD1wj7VZiBqCFc09+IFg9MLLyhNjTjMXGgD69z1yYN0t/d5ESS6ZIDZY6qt0U6yT2llygdfIP8x
lt465m29MyglqubNjsh1Utx5n+sDA0hoChEL2C1ZoEN1BJughsFBoik3BoMEo550nBndVoD+yl+9
a0JlD5mDOyWG753Cw0RvYrG/52IrplZ0baJJ4Go5NE/EX5s1ULECz3RxFhVeubVrle+FQdpXUyst
sm3I95vdI7F2dGP3q8XVdNfH9tmsrmNms1l+9BtSrU7ZWhiIjLUo1KOFm59YWgWRvOvulZqM5YH6
4PYO8qJU1Tr6uREP7XJ5aaJyQu06BfPAuLqnYNJpcSPfuK1/3zvni4FcUlFz+aCFnjbXmtt8cAod
SLeIkEDkRBI5VecrpPag2UrT1RnvJxdTLbu9i2HqvcRmWXO/4y/+/bjLdi1kDLbFXdSt5Dhs8tOO
f9gqokwCaDe2uECMgjdRoQtVh3pf1ybXGHpdIetMc5aRh+nk0zFUUvHbVkZWUOoYVNYqgU3/gD17
iafP8EuLQNWHuTZx6+Y9bw86Qvr0ogWu04rmwW8Nb+6sqsQohdMVxR4/QlLDWZHDWa2wv/CXjUt7
4mOvdOsqQi3YYkvyI6p3TVejWq7klILHEhkRQQLcjMRohfjZ7HRkOrd3L+46CBikTWMMtCAjYuAI
2B5mUcOev9JOqRuFRcwRsm03p3xndgxxvXIthRKDeeuHahL/QwicxJSHRYuqA31FUT6qex3WJ0mB
Ja5lV6H99txoIDG9tUlIp/dR9mDex22NNfMFTcJ9RsFS1CwvKmmjQs4eCzUzwpqmaHXS4owALunN
Y5SX8x8b1VDyabg8lB80r+aaCDc//XUdfmH9osH1XuYmfuwoy+fcS+CJCLzPKxSKweatiuuImkWm
jawRpH/4jxvjP39tY5yAP8qskFscjaAv7tmIRb33Cwh1lSbBZLCnRI7TeDpwNlWkt8GJKqLFLz5B
APJ5tln1vv83wSCqkO6xlJzSQqfg3uNX6RF5YEIcGyS4Dzp1iRdYGW7LnpzCqqTKQUYurhKEi6+W
WxyrpMGOd9/x9P++tgBXUjEd+ZJtuFGISVkgP9CS450UgbDTBZylNaaxPPWZchGvfaqL9HCrrQjC
kYwFv4kL/dEXq7pI3aN27fZFRZXT6E3iOIWVG6+SNZIcRHoBxo9IFooQEGYr4QbyKq+Wt9PuJJuk
93IsRg1P0p+H9hMGNLmBeQ8dGwUMbl609yX+xdFEN8tYiPBlQgt4BOdtmlA8Vt9dILrP6HMxfaJP
py2CB2vXZRgJPMiRXW3X1Mo1DSnbxyExc7q+TIKLSqCNEFGjzW5uEpzaV/Npe+WZ7SJOxb84O/XH
hs57tBeapjbZ8MmQ22JJQcvB5Nn1YkfsJToIrqMrxCqGDrh8en+06i4VcqQziKeuLp70IWhPGk/O
FKzPvPSVKp5UshcgyfBL0+zZ55XazmjswY3iG0xi4Umvom3miPqyURpFy5JVOx++DVEpvUqEhehM
V1JjgSXN8BSQbg8KQaq0xLXafC48GAWZLNJKJK5pcMT46BHS/6HzqKEP4btpYtRlwaSUDw2bYEEk
nwoC03g4RRIRRLi9C2OpsttDBxt0KUXTSuBA32ym4oUuqi78XadomBTpCbp3isSpil80FRaAuZGV
Lhgr5z61y8ZxepJTPiR2V4/zO2HiLU9WDE91jYzU0BxFbZr3otoalp2xSZMv/t/5sWDEkvVpI63K
7znbt0laQlypEpvw+HqDOaLHUPz+FwbGm30Ww9Ynm+6Nh301f+QJsXUZU+d8iWn4qe23BYxipceE
ZQNV6aLZ/vdioYinQV/oQ+LMBHXiZx4+/htdQFjPnzcPGQY3RVsjOhjenQYw7+n3FQDCOx2C5rlH
zt1DmtuD3beCNM0WStKSBcRjOZIjH+3evYI/SKh3CEn5nF7O9WPVs6ytRFncyX5gcrbhpnMDd0O0
kuk8pBpfeiTVOkTy0m5ivkRBl1OaZVVD3RmIh95RVh/VH3z6S/EkKLrHk/WV3jr482Yk2wUyHf0l
ZqYvSom2mu1FIC4gD2xDzpX/fcblXy+KN9j03w9F4wv9dZHSc/K3bjSMkdJH+9bLQae127myV0lG
8DEeiES8oZNXHrK17F2AvMb7+5q7/A4ui1Lfr1fPoDsHNsR2cePBXzcjFTALI1QvPzhuhLlItIuK
DT9+hx58JCLldgBLWQtEurX7JWLV4We6uKiPzpMjm7n20onwr9r2WsfT8WkL86Tudst43Sx8A9qy
Uo7U3G01aXv2cATW+wy0N/eyBFsVc7Ey8yrr1SWxNYUXYs2rr+iZt+tCEbwNIUy0DDWeML9w354h
CcFCRAlD3g7ku2wbayiSKDTlQbDelXhx7+u2dlEfzV0LfsFGmzq/kAKvNPv9ScBPZ+pK1cOkzMD+
zeTQJ/25TKujNLGPPsZYm5DgLbBmUGqj5YExFBVkZWmKdQRt6W6MdsdLqdiq0FJVsxfNOSEUQV5W
RxHV0LfMG6/+DXCwbjy2Mpc8B5gaavdjLe/wfcCpS2hXdjT8Zel0VcR7y9fdweB/1jMf1iROqoa/
I1aoVInX+Uo7Ke2A3TZLaYiXZGtLhW10plFoVm7x2tzYEYmJgOQQWuPTxfVmupXDl7d1aDAvhP9A
M48MpBmUC+HA2WRduQbxAfKswQOVyQMZIk786zjs/LXpe8m58DdwUDfxrKsUKatnN/M+KLemwerh
XeVReISISp/mXkebtn9dd+zEPP0ju+PcSsUFQeKHR48vWCtOZ6h7LWfGJTD4+e09CBGbslnqRydH
p3JL9HG4JDvcL7STnj2iW9gXIVP0cwkH7F8Ugbt/5LEZGZcDHt+t8dhFWDEda9WJRmQ4gi8UDTPZ
giXPWOK1FMpbuEH7mLbntjkkYe1564UYiP8hP5IHYmraXgqIutgdsWlw5+EsGDG4iie6vVAHVGb6
/e0gk6IACdvSYjW+f5DeBVdbamQQmQbeWOndIc4YbthkwT8ZHdXKrQlvp9iewdeBvgTIdhfjE/m3
kCkzPq3TRD4J7B8pxuPDypWd3l/PamPtcp2A39tR33V/0pv47aod3nbKP4RvgmE/+iQHF8H2N0JJ
ubj1iGsYB7D7s4q5coLURraa2pYeVctqZ3OAq4pKorNHVGHc1bhDRWizSZnysRcII6Chh24npLhB
k1m4ow5gBYWnvaZwX9WpZAO5N6Pn4hEmIv0G+iekSfmG+JizV2DQMPLKSTYhaikAi7D5lxVXhMHL
qgq6/lKSj3FZUidbwiYjE7D+ikWkYDhCzW0DPryUcGFWdLYnPWbw+DZP0ylUBgUI4G6AqEwMKkvK
qPZh/RvHCQsuJSi9dMcR3SuLrzzyddv70KcmXtTy/AfIr+c7ntTjHam0KCOEcKMj4CzD4rD2XWKx
0OoomYVsLQjVD3EnnAZv2wDyOgQipqtnseo0rP141VXXON30x4ShTAkIr7PGyFkIruf96k5AVY41
UJ+eB+q9MYZzsYqarczhr0i0bAqHJoWkCiD4sySS/22NzTCQJGCFiZPanZwhg9L4WSVRKRNGD1WI
YsMLcDsADPBnNY/z6XaVLrU0MSAEOdspozXPTfqO7pDZIExaQTF1tjFudsLho0mCIx8XtuXltKl3
rIvmln3GueXjW3LfKjIjLaZJHMDEFGyHX1cvlGvjhcY5G60v4QioHZ4Jo7HemLf5EbW7M3OQFPuC
o+Hr32f0yjQcj15nyXBxKr/im0tg7UFqU6IpXioEtqpXMLJt7EywMQcDYbK66cYFRt7GQt0+x+rb
8bJaL5KVAOAVivJ4oY+1R512XLVdACaYWYuf2RPnCiz3YzwaYjktprcs8ZuR3WXf1yFru0Az+yH+
iB9rQagxoVAZmif78Cwdk4ZeZFNV8Sj5SfjJVZGu7RpKEhgFAuTY90E5AnqPeo8pvZpBwGx+elVg
dWh6k6DDf4oOO453uvDhna/JX7HW0vxRJ4sZ4e4X/aBXHX3cwzDsvknHEQgECOjc60T/ptJPpclf
+U2K1VZTRq7MzMUZJhNLEv5ezclltYMoAnhrQks/6ZX8pYgLDnq8FgERniLlpuwkGaJyxVRMPYxS
uefOVVa4FxMDOfo3fTC6chVhd8fTxd0zOb9DaSsmIrHtFUH8qrxCLDbIw3TO+0yeTJgwni1ywMRQ
5AzPHUbBom0wU9RAZ3kJSa4klwo1E37+cnvmEW8vFmTBfS2F4w0HRPSsobG7RX8m9LmlDuM8YA3q
f9vER3Gm9rA+gsQb6NBG4Dai95/GRNd4q4EY8F54z2gh3oSsfmSnz/zMimhfywAufO/GUAr0GdCN
OI/w6uzYOGYB2jstvvUHbJ2Ba61hxNZXnBBYnJ0uw2pmRcymPlBM4A8+Zd6CrCxSF8801j33QNe6
swy6nOSnylM+BZKEQDCwjPjvhtIeHTnhdQNTZtlypMUXvxM0QRP/J1UX39h/OIIMIA5++ttq/y0M
/Elr8NrTfRAsGJXQ9T8wA+rbwsIpT428x6lWdDSDEX5Y0Zbhseb6oD0f4f4BVQmSqD6oYZoax2kG
2SOTZLHHON+iusy180UqRpGS/TfBlNXjofj2HX5I37UP9xTC1JXQrzyWIW6aagbEaWaW6X5Bx/Ny
Zz99g1U7U9HunI2R9koAENrKYAbPoa4+8Fke4CH0Kq94uJSZOeGE2CgbSiS6KGa4IzvLVC1O0Ond
ny+k3WE2jCxnyeT8KJFglepdZjmNQlyWwDAKESJRzCaEKAzRQSgN3WZzLBrPXyDekHqFGbI/Qy/W
EUjzFgnfKqpIsuPiGH8LfCP504b0fbUyIrnyJJuUitEscCbK51y4zomhv3do2euJNANnFVN4Ml7f
LMkojtAhrSmSJaV3Ij3V3VVbSmY3N/HmB+YbqZizn8iHChCyFD0K51CixCkiPRQFyDBvMJ/vmCJ1
yCIhS/l4k+04sJsZkHnP8yJ6uyxtvGpBsEeYtA4HrdpP6pQ3FKy6ZJcIoaVLNwLgnCOBvIhneU78
exJQJr1vZnWO+S88YVuLIPqaADySbiskavu8vcFYeYBZsMNFY/Y5xFCspKpWDkPt9kcRLxzyY5S5
ZBx65Uq6wT5Rz09NNbg+Vn/U2/CWpIkIgSeXEcUcGOcwhovG75GHpk/sRpnssMjYg9jBKlXtOlGk
t3T0+X3WMQoX2NF5BAHr7B9MXLriUdeotzIxdNj5vuA0cXUcwhBmG78hNAlwu+zC3jLfoO/YqJHd
zuQji2pcD8sxu24TIO5rG3eZ2IR81CrP46O43jNn1ZbUvg+Vaqvr+nvyfRph4p4wKMSfi4MdxPxI
JaDmMLiDoQmbDVSiL2gx3O8vD7rH6Y0miMrm2BvCJEi/yU/Up7J145lTRyN82351Z7AecafP8nHX
l5i7YVNuCZxKYpQJlsoPUjHeNbfrdAgRkBRennxgXr1ZVd0Q4IYgRujEV6yD17IEGYG6Uf1b2z6o
Rg8KIN6PK8saKjjXqBe6lw6kbmrYABQ73My2I6DLcTkVlDAQhsr4VHNBOWFU2cyqlPaMIYhxhcY6
BL/f8yIig2r1IT7FiGwwLhIrx+ZLAeOf7+6ucY7zyHG/YYkIOuFnpd9K20+FPOVO/Kp3n2nOHsGs
EJFKml8xRtGPDwvhrIiNWlWixwWs6iyxWmTO3ki08Swkdxad5l5N6OykKlp9W0K1NxwSEIbt0jSw
DnrBtfhjI0ypF07KkozhSjOjGFawenhHKX++b/VWVUyy05mD2rPnG+QYdBfDA3IM1fJulT3K/LEs
TKH3vmEfxsi7Xq+oQ8DeU2a5qH+Qi/xNt/9JKc3FgDz3k1LVriT2d8OZez4ByDUNHTbupZ12OAAF
kvhvteqSe4+QktSb3gYMZDhwMu5DYVPUhhhXN8UHvWrwEjkVZdxIPYlxQECgXPGqaOwqUSKprpjv
tldrX3NJI5S68ns9OSyz8oSxNKzvu+BCh/Rk1Jb3X2UjNrUqgTIsnXnqo8+K35YYECsm7AMMh93R
KilRm6IaqES2FWRfR9JLAEIIA19FX9sVw4NSi96VxQR3PefDVh/VrMnrPraBltn7yobvmSQHbYEO
tJSzMtt5JvAWGME2V3K6g2f33P+K/n/zpM/m68E04NFnWOGFVoNXOUWOI5k6fhfQhyZN+6GhDEuw
ilb/WTKZvutnOThcbJg0+my8PexyLdk9oVThSevT1X8I5X1gYO2vOAUIRQdevbyZhGNyAzHQnpu+
ENviSF8QvdGXfub8mVOdOuPT7NkLxYM1kLhptkxwri/3XZTvsMrcd73nrfjWKWaTavcAI/1earEw
5XFsYOlMrlaKVAotkOG7wXDjlczPaNgCRvprtQ/+CDT5TKDlMw441fC3wYch6EE9VfGYNRO+mXBw
xeYbcfEqFkSXwRgLKQE+x10SJ6NLiC/kSCqz/8eCO+d2RuJZlOi9w4q+XiWq8uKSFhff3WhnNdjv
XFOztbHgibd6m5FckCQVI0eCu0HO2jXqCXaimetxb1F8zqDjknHeEYzCG5m0sWRQK8wgBRFglSNF
Zd/YcQfU66XkWAxd6/99eJbDQJiD5z16K7FUg7+XG8TC2AzhsGSHnhhUc7tC5IVYdOfe7ZHeImwr
8msUvrE6WWGmU0y1+U8NQSBwKPRBB60JqYXavBuaAm5r9RwExlMGJi2aUTueZ1jbdPDkvZjxyy1L
G1eRpD/BfY+Zb3Svi8CZjaJR7PQmrDxoDXKQXmKubYKjm36cE5X3PyQLlmMfj/UuzHv8mTvAlgen
kS0ffExWmVzc+WHXF+caosEa5OxIIHO/h7uyOuzttYnlc6Vk7licQh4DdylcHzPWBypIDrtpHJKA
GqofsXQAC3jBtCJu9/qiqyJaGPenBMSfucULCc27tjLyQpW4K1Kvb+nmtgb6oGtuA8RwEGu/sumG
A2iVEAseDix8KwRjrvf+Y7ADCyjiQcOhD9QGqXnjc+vybQEqOA6GXWKUMwpnr66kEuNkn3A+RuRJ
AyYOuPxLmDoOiXT3c9fBGr34kabrckoFc8isX3sxIsbCqqWfs2seLZqV9WFii5Dbf4lcShHtIk10
2jXDrRZHNfswra01IH4NmSvWBaI9Kq+fWiAN6sgs2piy5LSxvt3hBhBtTuY0B2NjX5HWzkXLmSr6
k9cVj5EBd+t9e/uI2WcdBxwg8rnSU5TtfMBrxxUASYumeIQSaLDHvPZQopJIYM8D7iJASBzRLyXq
AGLgkBt7EvKhfDyh8lG9LDH/IsgDXkitnCs5FZaRCkE1LjpQHt3G0jvjTEtWc+h7hRGf4S+q4Rri
obi+AUkRWQMeih+3H4s0mBnlQ2rCsOSdeFBHTtiSUYtKfe3zi9Cm4IDS3XUDbGvq7kdxiQwWfFbE
YBgZa0nZDdlUU0lUc/GAkbv7haLI/kPSKHpBq++vQHJp+PYNnIstSbPhQrl3cMz7HnK23EQ4cCOa
e7QWdv7WqjeIKFxaZHIPFc0LvclFrweJi+w5vJb1d+GeJ7JzpUM3lrC/OOm3lFW/B9/S3pSn40o6
QZ5tsN4kkf3RKfszcuJmeiTXqnYolTyohgi4+Uc3fgO5TkfbMRYdwz1KOtxmFUdfEUnx9X1AiDip
+XQBSDdVvg5wL5epqbdZfy1OS2ojgALkhX7+yyznohGhx9Tr3q3kOFb2Hh7IrTuitD4IdOS0oMZ1
5sagA1XhZQsTTcPSn/ib6Y43sitT42CQRFdb9MSatjhAVyYR57O0ALkdWZ4b1iL+48CdmUA6xNpn
k4ReteIX0cCEAk6kKE65Q/+8+d+d6Vb4cbhbVCp0H0TjNqBon8i8+Dek9ciHaPcSnu0PPGSRBJ/W
f53wT7GlZDKas6btLxTgqEbCC6EGGWgFUILbMnm94r1huftC53TCabUpO56uZqVjj+8BAInWiqMY
Md8XMUMabUhK9T0WLbKBKBavjF7ZA/akYeZ43hGPR1EbWRDmc5ozwgIhRXhMz0oySY7zmJpReTuM
wxVOv+efF2ZONSzcYuQHFqtxJzvGgap/2xeZt+tEWgYQf14QycGfWjAllrp/BidO4WFVDagSjNPy
phx1uobQju3tioXviBNsHH0fq01/MhH4zQ0PgE5N5ZMoawH97VnlXuhIG7udbyayPlg1dVvo9eH4
pAuNZUk+jBkbdoM4dV6kMPzUiyQRm8bexkmtiVwFocLPeHMw/ICO95j9zsX92b9g7II8sI8EXAIF
WRM9scsqidd6t6TaCk6NcYs2To6tEwFgM+3qYnehgNSsxLEp04Giow9wF8s3/9x8xEroTTzOaKnl
shzkBdgcQakOKy3nI9vQTI46oj0aRt1we+xFDhFpyFNytxXWQhIzGLV3FqMcTxHyUPjwDmoT1cEG
v7M5uPjlGLWOFnKrblEYoF77vZCK9A+7yXQ5bvQQGdt+BtJTTdACbQ2edbb+mEPj9xUhMR9BRPQq
hODZVF36zHsmrjVTQ7onGWbHGcddywxT5qpVmQHHV83w0/5F1bxAQRPDHq/A0pYoZrhHrePsetEh
GiKQp39Kw6MSwQaYsyq1dhVaUY4x5QaNKCy6dyN4FZLuXdb5neap3IKFff5xxdqe8Wcw2J/eFOiU
yt6rtbKBtgRIYeMCQkVsMFCsjovao6+kstQqK5IIDSLFxKxX18X0JYPhP6zEzmStMpb2E2w1HwJe
QGcp0P7lFNtMmc3pEcqZg7okV14EHNXOuPGLh/RpcTBdLgfvKjSdrvFN+KqOvDWhvTLuVuo9AihX
dGFU00yg7+wiDSCmcS6LSOG6DnjsdkrffdqdxZkQxSitOH4Esy/9sHAFifeDaCd/n9Bje7NDVjKq
PS10joL/Ny8ai/u6xghpOEP8lnHqvorf6WkghfsCVDWDCIeerQd0PkD+nuAOatWTFOwKVYirSHPe
A9GvfZ8SC4Xc7wwvbFZpYE/MZdsnRf+VKFlIjx+sKb2b1PfYkgm3RH4lClEPGcIb6qkZ0DuGBGYm
zhOThKjXfm7JLbAPS0mRTOrJaYtkS/hmzrCVCcY0wu4rDepQxPQRs7QqkeSZC/YvhVLW3cDfzGth
XQw51Kwh+jfotjuBExDwNVD3RYk9JGQ3Fkr3lEDgZiIRlB60q5L3Ry8iD+nwQqzkQDOcfaZUsSVR
PF/7gFkWQYwu6doSFV6GV+PstJ4JeSAbEID00+2dGaR3+iPQ7W8/qWiGbAhgY0zw7ZhZ4WvHhuta
npERtWxDsg7rh5gbtlk3TnKIqivzrv4eywZ9aVKrbC5qKionNBd8MUml45uinqriu1nLBiUvG91W
pPpyvVJfc8ZKOj9mQvpKUnlIV6gbG4Ny/5uC/gJfWYqY//NskO/4AIkoLcRiQWKsB4nZ6QDXaHap
2NX/JVKy4x3GqgdFNE0xTYYCZ4Qv/L7YgajP5ig2YEW9zJy3GzIb5Ypaw868oIBiCZytJAUdad+8
VuDEz6UPv9O7x1Wf1nBQCGjgcc4tFN31Zuh4I46n3eLKpLUzd3KWct/ATTchpoCECYqxgAKUlBv3
JvUCYHBIhmnnmxvW2h92+oE/bTdBeFtbZnnVaOE2vihvUh4JVepurz9b2tPW8SLQvcg+7KGIhv5D
iXUCZQrb8IyVv2oEqsyKlsnqO5/fGLpLHgq7sCAx8Gq7tTigPnc+rXRjJSUBdwI6JMmIVpiApZ6G
wjJozoa6RKlmJMdw2qf3JqvJUzEuPUjitWaV0VKltAcvTfNEayuwp+D+zW2LJbXXfu3t5akuG0BH
g7GradMaHcMA8Jlo6UW52nywmKsfnkSw3hlHvblQVL4e3mobqSzL3d1Y9agCYEcsHinILSPyUMhX
gCOPkbOB899vKw5+mCpN1fbo5LO2vGO3J2XMHttj7qEj6cTu+kuaTdh8SVRrqhw4VNKVcb8NwNev
djfA3I06OSvNudKpkWRk4x9Ty27ukSNhPNmWOgD2CfRUd+KfFdo5FqGP9RSCJUHieHifaYi4MQIq
NTAL0NYLfBJ9ELA2croPVftIYvbWAkDpCM3tS/+GC97lKglYZAcwAnUgLlpeQhHKXWs/lUyJ80HD
tM25SOgYNjAEaueCbrqe0X5FQ4oShDFctt/RPjcgFHvIbynfSgK2tac5e3Cswvsg9WCL/9AR7S3L
39zgEennxOFJblNk0yhVn+Qc69X6L0FX52/a9SPYL1Zf+kuwMKJkPKxMpzZsGhiMVW5UVArZcdW4
3+8HrL3xxV0pOdzgHy0wonj9urmwIKzLRGqAbame3aMT9cS4eXiGctZjT1RT0h5wRXQsQ+5lTyhA
3MRp0mTf9YySI37tNxMA8KLY0Q7N+apwf1lUw9/iHoMXr0WtgnQqWLd0BauaQeIpm964j/4+TF7b
1AcsntvHQbKQU5KKE7qSSMU5Kr2B/VtfOctvWnRDwG/nMjMlM4X5FNuvtmAr26+cLhKHQlOiywcz
Hg9RZahH73dUhtpMYPEDO7LmAtjO56MD3JlTS8eeXcU7ot2BsIJfbi3mJP+a41hDj1lzRKo7MO6e
OKBOLL0wesCqGke+YY+Ujo1eCp8WDveyC4qRyv8r3UpN50B1Anx/dxsF8CVdKAGAggvUdEzNCvui
Iyfk9AGULg4yz7/qY/IcI6hsffkcENP4YSPfPh++ehWyBi2RCxfCVF3N2jyfvHFf+YZN8qrlBr1r
U6+dUqwtL+1Kd+H4ETNwBuv5J/ON0SOiJGciwm2J6QlOtJELYZ19FWfeiL0jI7lsrIaOAALdFCYF
xUOnzlD4zbjPVCJaldggW+BydU3vPC8oxoELPlKdDMeDNdG4ttiBy270gdmq6ufCrgPnFUwgPMbB
vrzhDof/di8Egob+t6neGuYogDPe4jYn4Nz/DkzKiO3UU8Gc9y3t7ftxtBTYynM7gPUlU7H0ubIl
kyVik7p8ZQYJe1Y8L0bNUn9SgYj+2QDoUBc0thw8wpl1S1WSbrdJFoYo2Snn8j92wsxEXkRFvy64
g8l/F1pK3xyucUoylwVdHgHy1kZemoS+aBeZlZKTweoSRBFyFk3g7L8Fo6bT4YYKTpYp7vFHedzR
GlekD+KnQ99dlqavNaNx2/x587/KtA2ono9HBYjhyQdmxFmMUx0hXR3CuMDzsp9Ijs7SwbAuev+F
IlaOwjaYzI9wMSLVSWxVitW07cHzuO27UmCt7foTeL2D8PccxmcaEGWRDeeQASQpOHZdPgGjSHEI
hs4+dVoCvhe9iO66e+7ba+QAZ+Jinm4BurcsknAIHbdtAmTw6pDTUP/8V+eTB1M428LSAMdsDuJr
qAgn7KgWQ15ZUFFPKg1erU7nJ0RkcVGdvy6NseE76I8SJQetuTwn9D45UxevrzNTyl3C6492R7D8
D9F8UhjwV8GTkCU/AvOqauDbjWEJy2rBfwQQM6XR5Bo4qpFwnl1EURhh20gjS7afxFk1kuCThuqV
IRfl1wkL5vKmlCNuVuSRat8zRKYTK4CTKcH6LwJtqdSNvmXQsxn6RaCny7mQvUOrPUSwyehyN5OW
ehDKh5nU3QBpCTJeG0cYrWyVKpatkvMzPSzPpenDQE+oSLEp8A3Y3O13nK5TXWCg/C2QUsHS2IAZ
3JTP7jlkROy8mInY1XxbdMpd/vhzYOMfTcQaTCHesMzaMNJS9Et3F8nyl8ATior6M/Flv4rCWEx8
EZNIbHoU9hU2uYLmVQKj7i/wFmEcrXuCbMltKZYLOXmLwOlCCw6l00gDc7Drz3P0oVTzCUhLmsH0
5afpEpyDSxkKmoPcqGv4ObPFTJt9SY4KJFYE0LwVgOLNSZyx4GGn/brHXr0b04k1fjAV0P7kazJs
9xhllHpS60b44K0TBmfMTsfttEZ4WnXJZhP8Nda8CfmOYcXnXPzDqM3jIUUtYHwdGfTijhQm7PqR
zwdG583BtbtY+o0Kop05SA0dPp+gX3wTGTbwdoP6gERzSdzSnJIQi0IDldmljG8SfnAdwFIfxKUg
GM11Bi+jmqMdn0r9RKPGzVs1BKmf5K0urnfbJTZht0jP3XEztNc8wiZH0PocHvbgzSqErMbQypOM
hGLvf7rypeY46jNpUnpwYKZH+iUPdlwVURAo3KXD6g2ROxkkKXor421cXmbozsRYGoanxKEhanSR
OrVIE7e29OD7Yp2/6qu5q/xaUxqar0UIF20iARbelhOFiwBbFaLPsLuFDmPKkY4W9dbwlwBy75kx
1QSqq211F9up/bShYOXFCpZSomAcXiVJu0CKtRjrJ9alLXlTfGfjpDoO4svMKlihyXIp94292I/b
8e22oU5qbeAfSJzrOWlJrsHa+6fpJWYHJYwPtUz8PV0h3DkDxj2JaWgH9huCmHzT7RbhSo7Jyagq
ho8HRO/nhxKqxfbAok+dNqYcUVTAHkhNJUa/LS9UCBj4omBRLp391oSvDOyitpuYR0VMDolHE2y6
LycWBEm98764VWubVP47rqSEPlSEbns+nc43PJSyUkox3Zk813gM9M/qDZLDF1cPqgnHKWuXZtzE
gPPWDbVHHxvYsUaziEZMukkmw+7oP2HvNyt5U14M2CIaV+QrqiJ0uBeuRsACvv2OTaEdXO3kggz2
UI8wcljKhtPVTLPzVnvTsUF/dsDFIObk28gcJU9IWzw6SibXk1eKidzz1rohvWbCnA8sKVLUaN8C
jmAH2qP67rtRH+qKws/3PtaMYFoTLWhbFWPRJuTkD/SgZPD+O448599f/OAkJMGQXNwiXqPuoRBY
k97Mfn2fjEVYjTau6+Gm8UbBsVSuMkveMI2q2v3EAmTCGT6OYS7eKZj2Tu9H6p7SqSsd5wcO6f67
goeTXiLl+0p5woT4WaXlv/1ALq01QJcFC8PlU8cx5q/IfZrsdh+4rxBvMz8QuQzUB91kbrrUjks2
B9cDQAtJyTg1Xst+Ulk5SqGL4ox0SejXpbij26/VzyzHZAc9sei3i9zHIVwKDgFo3iSAOny3khpB
Mm4bY0NtlbUpTX9ODT9IM9uewG56bsIowm0Xwb9ZitoWfhgKqNXv775QAcUQqyaydVh8VIiaAp8n
kgBZ9LFHE15n04VnqLw5ct39VnXmXGLpCWfjAZ4TCsEanQILUjByrxEikW5jOe89odip5RwLsQI5
7ZUP9/nQ+Z8KL50ZCABw1CVk+Z7KXy7xgVUxdU4IOSPhiJcS7LLZMi1IDIS4dplNEjceE5Bfq1+H
Dol4Osby9V0zOY2+2AyxEOEEbZpeglU/9gP1tKpDaXwMcRi1odqcq9TJlwj4c9qPZwYk1u581w5H
1YJY3YFHgzXA+wMZHt9cuaBhoKdj/EKXSDbWhPomXs8hrP31QvWMdLr15t/cPYaBRT4I5zZLFher
JjXCxo85VXTyFxupbATySg1qkQth2LWqatlTZ7UZJS50Pw1J29N2Zn/OybZMELCoyf3ZFhxhOESl
WGYrpzUCCzyVRWrD1dv2QSQUb8A0pI+wXPhgwTTNnjdhemKbR6TTEpUpcbqtnQYRCAphg1vPIknf
IznUZpdKqYSvE1VBtwUPm/CMH7PECWnv70iTve4uRdcJIwWwwgVB0gVDDIZ1xPXZQQxYoV3zIIDH
Jm1M4CoTXjv8XVQW3RQYkGH5w8k6wOhhxdYXisBtcW3K5Y3z0UW2JXbJj+chJ0JRj0CoK4ASOjOC
Vz6Z+PzHtnkk121shVscQuBbhk7vcJUBQLZhcKgWHcZsZBds0z5O7Vi76MfjUMmJf4AqC9C6asm0
jLl4ZoGIHkDrPQ2bCOSOljDXP+nyJp7kzCTpLHcLr4vFbkybFM8m/2r7g/cO/FqQomJqUumzIMBp
kMjX7UwBxiPRrM4mxllFc+viywtkDkcMcsYLWNMIzXcdJaorPknrMS1CLO5+QeEuE4532lNmdkPD
TpjVY9undYHgztx9m/AW8mg8TZRjjXAreuoIX073SDfo8NC24y2VdnQk92a/deoYbNR6eYBes5Qv
6zH1+DO2sPKvcI84VMFHFWOueuKLRLfAX63tVSaxOD5TDFLbcGAdNABB4+MXWVs6a58WU4jQq3hC
I7jcj3fAF1bghF5vyKTVKQe1Wa+IVP8k/p9Mp6tXsaRy1HVJHCYCl5KcHDrIFdB2ht69gxX5vptc
fFEpOdR4SPSs7yGBLO5/rGhLn8YjMYPSJiENtjBDxo+f7/eNF4iFxmqdFquU8ntEDj0vdGA78SiE
LIT2f/X+CuphAVzP7ylMe/FaOGmZ0Wf9o47ZRV+8CN8IIUPtDqcW+0LVkQxXaibs8iJlU0HqvnyX
Ed4R7IkXFNrpisFRX040kv52b1u2iN5WVVGkNGFNT6t+OEVMoo1LLTQ19BK2QM0S2jvLeZBKi8UI
NjUV98r0Eu8LDS0X2rpDowt2Ook4QCs0IkbNduAZl5tfmBqla3KpxmBupGXTv7p66pr40CfEAqJn
9Ye7qYfws5pdR3GRJZ5w5ADm4cfn2s64tAgvEgrzu4EgDOw0T/mjHuKlcPYqKBMXI3UZwWjkwZjh
DyQtOiXHfPxIIEKhcefbtZ5k2oDNUHgCln9cjU/8dtJC9YYWb1MiIfvep1UjZeMKcXSl4i6yhfbm
TzG+QY2lWmQFjQ1geYmxpS1CcIJGBW1Taojz1r5SLI/Jf1NFtY0ZCMuC54oJWvu9zjNJWREo4Akd
NCJHd3b3VVKb5kw075bFsyceMpXRx4IHiQ9NdDqevgEYpZHuP4SaCP21s0Ag/S/JF9U24ahsVpS5
D+H1A4L6xrFgyp2IFCrCNCpXoR+l+pF2WZc8fDMnuQAeKcec/SntDKG8BzBwLcB6FhUOOs//CYwi
2LNEbJRB1PMmjqFl2bj6sFyOB4S+/VAwlZXio0TF5iit0tNaLsrFaVS0k/beJIbPMh9OLpdrpwzm
rtgCKQVnxlubpcJ+VclQH4aGnnf2pvZ9JThOATfOSsjOdLbBS5ApX99Nbu0JGNSMPAcSTrtxUlNG
1oPR+DXOL5UfokZXWDN8U+biwM3gFXZ64P7Ptd7ZxGkSgcZIYkN+gn1SKfS+40P7IATu093qBfN4
Zf+lKru/tM0cHX+bZLa1Jvyl55lHtdCv7+xyafPsowTLwyjJFb66IP8xGgqDi7fph3btO8eJaIpD
7wFo29tRCk+MkDXAE9+9MoBIPl42v1RpUgvlxV4NA3Q8l/bazAA/yvlr5P2Ppv5ZCpd2Jq2hMqIj
YrcYSnnq/Ms02fiVVkNMGarbNjeu8X0ejERRsFqMYU7bFELSZjEKBxNUZb+yk/OUrM+w0hJjXBUS
/wfqIT3yUKPr+kYOteJwNpMlABUcvRzCQslZG0xQaSRq0ZS3E6fKBLHjKyp+OLxRLrH38/HB0EQ8
v3e50sojuaEZfV6FCZ7EllCw2HLLXwCZoUL29HwUelg4SXs5yqJpBXNtwGjkmkRHmeKiyvKKfttd
LmTCVGmZQ98+vMsankXskH7VSaD8bUeJDY5EBr29hHQFkouDTGpCXFe3R/vH5hrzaoTjzXmVJHnh
n5joG62WrSMe2dD1OXzoe+k6PPQ5PAYzoFks+WPZ1FycUhdWLaMNj8cv/6WuhrjHo4MU8OoyqDEo
KqaBso30QvMhVXuMC5P95VbUdzMdV3TItU83CVB0hHsSTzLnNKRBxgv30+qa7jWFjIyRUUEsL7JR
u7t6xavy5eHuHNL9+r8yJENvbkaNtUf7F8ZCXhBOBq5kSUWorR0v6bLfgm5K8vBfwkBUuD7tCxgl
M5xMjpwN6XvL/BpJlAR0wBnKeOLUUpmqPPfx6+5bzndJjLNxkKMzlRCm5eGwnQqVNGyKS4ezyGvG
y67Z4b9p2x1VznGwvmtvIBc04l42EI743DY9T95/s8Ds8qTLemlcJSss//MnVM5v/3WhnZWBBz+x
2tkRtRyrnztmd5rC+qbasE2xri0nzPB0NemZ7zNuSVx05cwFsB3PMNG/qzhOpGf4HOqI1TocZO0i
BSFR3zh2/ZAtBvPycEPTSKQfYRWwLUVNTl7jOpX1n1LHtNI/LJY+9TesyZEXF9S9F+Vv/g/Zp1xj
fnRg2zeGz7HRETsi5CdiCsk9hToJp1kg1excHl2eiU2RTbeRNEbMuuymtUmzEy4fASSFG669m2yZ
/RlABj2+dh+UM6UuC7BMJFecel9uu3xqowGb8u68Q9eHJSsPQb3wZa2BIwQMwr1lqxeSV/rdv3l0
ys305rjXR6upNCTVTX/KeCvTh3WUVYiUnQRV3bsdDWT4IhX5RmTej1Vp1gW95tvvsN1FuhrWkgta
IK1kpU8eu8tWGOtGLUhljyASraQ/hd+Y3UWIuA76zwm7PlSe7qF8WC32L+wpzBS0PSK6TgXnqRRp
tTJyOm90naHscO6b9NeiHQzwDGoed6UYrOA0eM73vKSxyVH7eRHdRM7etpA0IfJU6y9kWIr08Ks8
/gNEpJL7x+F/r4x6GDImLy8v/xSVyhv2roETdrR8KmnvU/pkuZzEAuqc0T9t3/U9zmkVXc/7VH9o
fSgNDwvrEap0IZY1+0pz5DIV8RQ7ryLNp7GjYGhaTkrGHXIRq89XCsvfnxyPj2hH+aS/XJFsDXlq
Ntk7gT9927oHP0Brl5rilYVgUVrbV1vcaZ/EvHQxienEk9VbvqmOnzk9kLo8oyKQA8ffQGsbE3tU
y/PynPZDNChVKj5EkesvTv4+xnPuXeyYeWMeX/S1FPlbiQPXaizq/PllhBDfUVTy+7jvJC+hUTaE
dT/pVnpYtvPB6JfW51SlsBLt1RHE0cafWSMIA1kd7IT8AveF8BVY33JBesEOUSOTlS7KAnEnkPfB
MziaOk7mjw7thiJmxE9JVJIhIk0rMPi0R2XmQ6hf3OP5B351y4fbpdwJ1NUjucKPM//OmjvX2ezt
p/e8KCspyqGVqmEIumZGxNYPMd7BV+tMJa2Lt8Fk1n6ZrZVIx4D/d8BXmohdkffFfFutEJGsZOVu
9/llIgbPmsPCa+tUS75I5YvdjbL2eAwlbhQ9C8wzETY4uiCreuehpYCmA+sVwBfD0DuQx0BLl2zN
XCyarJBx7R7nwAOVupoQXX3Xjd/cBfg4GS2fPONhd2ubflBomFqi5OjDyqWsfMN1Kf0M2ZEmW69a
GC8m0jRnh8mMwajHSS/nc9JwTX9bH0L+MUj2reg0jMz8epJpIbNTJMBSA/3dsKdZjnPXBCwgIPHe
Z6FCMqRdTP0qV1AwJNLr4SzxBsOLO+nrdWCJ8zkRq7z+C2F4H7ryARUnyhl0R5Q9yH4jvlUfgmZg
i2Tz0UsM3MgROEUf4Rzs51yHvBWttI7k0Sy/30VXpBfeDns+L8dBUaMao3dOgKPYiSCoK/jmuQoe
6qykaNI2zIBybtLAaSLP/oaiRVWOrJ2ewdEsLyZinJg8nqVprLaXvT7hXKKdDJuD9wdFNsZyRIka
l7h28l6fsLXpZpvOG90PyWjnD7qjj2eoy2teb5LlJoMRlgU3uuPhf6fiFMM7I1ciDEsyEuPpAEKo
WBJjeUz/MpX85nQWJkaadgFUQ7s+cJ0GteNUF1O2tz79C3CETGj6ud6SbxXaoo2ZvMUmRwDoBxr1
WDjQsADYUXRK20j6PVwNN+QP6LIPTya0P2765VOSineLI+0XWK60WLNEJ7iJfTDiyzzM6pCHZPC4
TqzHQdN3AEIZHJNpnMLpZDSCWCuwjDfMKFqIW0C4YUmY73bbiXSe4eahQa1IbW51j7x9TAPzZ3iB
TgY+6G9SPNHznIgqO3pVkJ2eRWGQHSev6MaLXIM1j2nT0T5RrPO3JRSXCiFb/Dnkk0pZoZoxloWB
cY1GBTqDwTsJbcMrb7PfDb7Ce3yNYmPpt9bf/eX05kdkQy5QX3UifOY0y6fnSwFV03O+MvUTBoiG
FnOYZ0TU2jNJDes60TA1uu/T24TzYH6ykZkJSIVhOCMwHIwX7GyUvzCWF2bDlUOa2mCnEhnwbXaL
nkvGWwf9nnKuPWKzxCuRqZYlZHqHzR9NqtfYFbLxCke8WOKkomAeQYsRA52w1wwBJHrg9G7zLP4s
cdUZbia1oCi3SBGLNWSqZWM8J7yH5f58hYZv4FCokhVvARc7AaNxvl4ZIaUF4MHXQb4SJExqTgWm
k0kwZQak9YZ4CCKOzWdAosnSEw6tY5BBoQGvH6R5V8qjKSJhu52wyLpP5VSeV6WqqKV9uJXV6QnB
V5lkc3oYkY3aZczKZF/35p6rdVwFdkKPyUG/p3ge2uCvx+h9O3yi1n9ZkfL6THjISPoWymInSerN
ltf+Brr4HnHtYhxCeU89l88dbG6i4n6LHEKzlk5H3QCXEEdK0/IxnixX/w5tjzyXLLQR79GZesHC
BtJM3fkVwqEVH8RgX0go/oC6IvTNrXP1w9+2xBxXT849ksD7c0rvu8TkwYS4iHsqU8VY9fap4gNJ
9CCjUx5jVBppuKoobhi1smp8HXIlN64PHecaBC+wSiJ7s7n/blTF8xuvRigKi5R4QgdskDI6dyA1
Whqk2Qnx7+GSexMN9cBirvb9DxFob2BS6Kc+sNEgF4O5y3WS/pzCEgMBqaoe2XHvCTIfFxZlIx6a
mMD+lvj2sUVmGSLgK1IuW6mbXAKZzA/kLNDMTcijhm6PaJeYMZBF3DD6uwTkLUXOnKndtDt4gCbk
jY7erwB6hoFxbCPg+rtD4JLPS44V0nPAjGFTYCVFPkM5evCRqRx4kEhRgk2jQTEUlMjzZKNbmr/N
tG9NFy2NE9F06P84iLHO3mOd5q0AsR9EoTWOTd7Lm+TMW38Fw4gR6o7Uw72nJM3kT51+ZlGLnGI8
HQ3JvV50qk2m/PjWsqA6zkZQx0JQLvMnfBiKG20r5RXMuBKbT15YwJ+GX+Kaq3pkwqNMueSEsR3S
HU57ViMnV3Ax09DxHuY/7Va0pSmfTTVQ0L9P06U6+mJ3RXEtihrG/U8f1s/AT0vCgvhDG44llCfs
kXw/QRdXxRAs5HkC3Ib6w9EKSI0GULwZnkqrdBcIthkTciU2syxSmGqURqdDsJB4N4fVyLbhQD0p
T/GfdLzYLql0Uktit5pL6FW5cURYKEvl4q8lmyY298N9XCDqpzwIjMxuw5a+Y4Z5whBrLGA3Ibpz
a+xyEg1Hc9d9G2K6BKGVM1/9sjjCUdj5XDiIgGktT1fgqvnk2SqIo9thZtQfX8R98csIM/Mfbyhd
XyB4FQAgXG9w1u7U53yAcQx8MqQ0OoEnwsToooRP6VkOoAA+wua9BzCtU49Y/GCyzRFAivGwYbv0
nigzzgBQXVMYZD0UHfjtd9pLBvWo0WnnK3nvrwD3r0LJXjzRclrFkPr6IS6UWTylydbNUzmwfxfL
pASkEbY9vY3Hi0P4S6qlhY0XK+OTRa29Utx2A9WAXH0dXf08hLEXySX7mszwntXArphrQx3zD0Re
1D24c5QbDhUtHe613V2Y55WNgsnNBFJF5bTwe58RHMzgYRe7uij9RKv/F5egA6ji2gFhWTA9KiJV
zsRKLjbMzqSepVJ6cuHtQOR4cs+swdfCMbuzfe7LDmcA4QhGlXoRinkGcnPTfHYVdtdnbQ2PlXzk
uSSAMrnoW/Dlvh2TNExkCxWJ8jIWCVRZ7nleFCy+XcwDqj7YhtVpd8I7nyNOauW8ettfq2hxsOo+
H0EJayRk+8VXeGh51SGHILWlISWVNz41KTPqvWVwYSLNHSYdHXJ+sQIaYXXhHAq4Cq+kJ+sTc3wr
2VPn8m7K9jcP/Mc711FxuQdzOVUQ05Hy/HeWWdC7UA08/p8sI2f4hcOw98bEC6D3tPgcnf6+zYEq
uq2eZegOpznFxO04UhkFJNQ5tn6c/2lBZ/cDsffdyh4Dc/k71sBpjxVGr/lsyX0N7V03oStaPfGl
R09edykYWmppSfTZH1TosVMETPP8acFlO/z/WoWB6l/ZwlKM+wNa9VKBhe7t1IrEnqXYfBrM91KQ
IM7HIn3jkR2B3Vns+WFkd5kLQv4gfvAWeTlaUn8FcVSO9GKsX3X1VOM1JVc6Jd5KDU3UiObKCfCj
S8nLG7jRsIHzebUVksxVJV/TPlCcb1395MiWYy7lZGDbnGKAT4+ycJdQJu4ItaUTVtw9HoG2gudq
Uc2iKdSdbmJMvSITq6U10KP2hn+PfzpHbjODSBNM8xIWQ7oBFnsVg4uMSqK6E5M84BP8jipnrErm
Ejn+yBqLv2xiQJjT7T86TpHjYVSwAbyNaxztImNk8UyjPM0t0dFj9Y5TBW1S2fpDnHhQHXq3rBXz
bjYxuUYSXPO/UTSmCG8XLmDPV1p2QTJCtDN6S9obT9loPsSIY87jun2EwEPHl6bc1sy/5IHrb50R
agiE86bJl5hVyddgq/z7lAf0FSiGSBHruTjNs5Gsz0pV8fwAifvbiGEIvuhHag7nBjI3pNb1Qoys
1r5TRLe1LAjWTnX/rgcBUVSfh1dnXfOxkMR8BAh2trqSIsSq8hEubNG18W7qyG0xBN474DGc6l/A
SpMZPBVqz3CuMAtgnp+4tJHh1aOCM5nCFaZcxRP/9/9f28N8rmrfebZLrN0jnRcBi0K6QGuhXlwc
nFTIoOfTKIZ0JQI2udC0G4hKdLmdV1gYURKP2ojzUFry96Wqt0Ru94ae4PeaIeI5B3k6B0oAeQFq
hi6lkAPZykzAuMkByrGFZOkIoNqxx3Ffdiyn+lXPqPYYyF627YRKCVvPtxrUXKZvSZO9W48u6wLq
ztstCWjDWm6O37FQEcGUGDZZdUB0CDU4rl+ovXAPtYDbU3ERtF9VCBZDka+fS4sSmpcm1T/0Mi9T
iiR7d2NbDkdAVAjbGgFKW1wIEnXSPdrALCAtv/PxV5nuuSXBz+zUzDw/MSza+iPg4BW60gfALXSM
CNAGqf5asG3wEe7Hm8M0fb5GULbtI0YUYSIw07LQfi1cbac9qmEH3QVWXUkQCnDXUTTignbSFJWP
hBdtCDG5AaVociKsZmlDqt0Qr0iqxJdBRoW1ZnLakE6nVhq2ZiUeFEtZFz536Wp0qwGIhzGM3Jzy
4TwxY6I4Pnrg2f4noE7+7u8djhHEKINvQ3MPXDc3VVi8mLJfnofH/Cdqwv52/sgVB4+vLHE7apPZ
fKxQRaeVmuUNar4fctbOioHJB32Ftk+rRhFT2dsZ3YZWEbT5In0/cy0BQDpFLcKRBcJZ76ntROEg
KimYdVo3jEXC3He0ARsdU2c4Hk1vXKc6lBtHHbDEfYEJN00QzwdZMKOmWSft9OI8r1m8z8zT8crc
vebrfCf6zFu9ISi/VDuTgxB0oBZWAfmA+c2LOgN3Xuc4N+uSIwY7EGg9gruV3wYZF4phKln/c/O6
tmhGkHxwqGRFVGL8YQp9Lx5eqctfx4HGhDkOMlZtaL/fs2m/qxJnYYc7T0ONvI4/hlGaO9JtdOcR
3GuU5iLiSDJWw2mdyrv7iSOQtYmFrqscW82UuiMqY9RKcj2OUQPDkCWd49vsq0iXxo2canMaQF8m
9kaWBa4Y4eayOtrSNCGUXfX9ttfPJ0OcK8+n6LBt4QZuODmtIo/7OwJszblBCTYTvPYD7YDanxEL
VTRe9OkZtGzc7GO/wHp0xcbxO4b1O63Q2miKIciSv5lvMOX7GI3QuIwit1ASAIaKv0BWXvzNuMT1
nZb6kfZGhurZBrpons/fFHKqMVbllcgVr5zcAgB2qcnk2QarYpG2Wq6WctG6bw+QTCdXzjHCjuAd
xSM05M2b6VaWxpkMEfvJ74O+mD3w3q87QhTRf84pmZR/uoD7ie2Awbz1thQbb6ADZVpggv206bJ+
n4BbsL41YCCTSEmVpm6uFGv+7uDjcBU8OIjWaypuOXV6VsHw0p/ZAz2m6u11/3DYYaTeHW7AmiqK
Zs8h+8NMrQYcK4zR5MNE/56nIDbny2640/0yDrcsQmp+xNMONUmngEgjpK1oWLYUn2Mn7Or99oHq
u6FAzNOc+8SUifn3OAl3vMk0vMV5t2WtXILYlvg5iWW2bAJvCWSh0QaKm9PycCKURWLDdkS6PGc+
0iF7B6jkO5iqyHPb+zlrTNODSewULWx20iUum2Ug6dg41VecZTVoho9j8bpR9go7MVN+7SIb7XoU
j9I7idEZ/qT39DijxcT0MmEktxkLkB4ViQZpAyO1DOQDO8fQz0M4Z1SRnysnEjuyzRdh1D0tzJmK
IcUWRV3pOTu+Q/zEko3cQokfaa1AlfE9A/pWuOWrMHyY3q1dMA9oFSt4pn89HupghsAtAV/D7fPc
pNAMorwNQ2v/FWaBQnUMnJopL833lkOQ8wy1p6KE3TOVx0dRtJdRZeb4eP0ChvoJRuBJstmqhjKL
I2LoJuVqUBtpHkIOmUEHtmwV45ojHYeI2fltTKBSEXgsmeXMb7gPi270I150r+C6kKccZ/N8svTX
yUCm7PhjCtT4F897W+wlP2ABi1AkDDufYGNK5WgHqwh8jqSCAwPNuGD8HYy08y88sII9f54YhKg3
gk5iVGVM3GrHrwZcuTF2cN4hvyqxpyW1pdmC3ap5sLE84ZEXrkUPOIcJRcw/26zm7fWXRYvaW1yu
iZIR4Hh382pW7rHTWriFkqaa9rDOD/YP+g146c7lfpY1JmQOyPJsRICiaZu1fgeDRp2nBiaAKxqj
6jlD4LR8jwMjIi93KAY7qu+7R1YxFMZo97K2IKdsNkiLVBOBNDcDG+Y4kUxy97MuglizgKQnrp1a
FJw2PsX7L8TLYMoSwe62rgaZDTdWwtrMq7tfuErEjjV9DPi8t1YRavEzuZvMbilu+f75J/+TuOhU
CDV8KONQpb2EMhvpsVMwFRyYVxjWfakeDp8nsMXvPC6MVzSQDE4k284bmzTU0BptVyuWpsQ1f+Nu
ti7s/qPHB7IfkC6nm2Rx4CLED+j/f9nyaZtsk/CRd1So57TzdF03QGxlWsPqp1Htgj3+V2ujVhYb
QTU89ok7pYmhVzDDSxx0uEKRAhorYUSTevU7RDQPxWISKyqcSVUpL5jmFUC+ii5LhfcsWjx5zmqu
F5xvqbY8lCgJpBtE3WU7GVtqvvW6AAzmyEVRO5NPhBqceoqADnb7Ch3l0zIoP4SAWGltTOgleJ1z
vhs6IDFFhoVBCh4QT2mTWyYR3ZcnUk+VQviGNGh3vCMAXVS3++Te74k/2uM1XeA0YLy04AGFU28O
w4PhZJcVlQjkOZ6kQ22HiqNNL8YYV3zEzxeRHRvhkNp7xvOAB2zGTH+bDS20WJUbPuyM4V2CWoHp
jl/P+KbXof18mJeSMuWtZI1t/BES5pPbyZJy75OLfTze36RTylQpG9CMLLn1COaGRptreNJYpy3A
nrQrJqkSzpBjcHPJ818XtMuEoAQRHYxv8gqdykmNN7gi8UM95slle9xWK7ntgfydeuQbYLarPhzA
+it+v9giUJPfLLc0pb2ddRSbHLjyPLVF+SaJkPEF6vq/n15V08zwSjJTgPZnXUs4xKOvP4RuiWNP
+Y/mZljC1/bkc0hPCaQEkmR9mjyPGQQxmur7y+SKpRdZxUMB4VhUR2BswApz1eDNr3lEugl8KX0c
+9m4YQkdlt5+nX52EaS8NIPfL1aKIz/iokEU5QSEI/i061wuf4GXUJLXGyHLIJY0+8xiZkYlrqO0
aczibw+ulKqeGiYOMIaUP2zcwgQdg3nj3SWQpwavNm3SPV0h4WubeQO6GnmKrLoqlCse9E/SH4+y
gg2iH6zPo+Rc2eiZHGBYBgF200WKgcO+liLTjxWJN8tDl0rDzB8vXO57EQtkBeBmyVLt5DFq0bMV
1IhX0RzEsQbW4ypPK9U19Et7rOjxSXD7Dm12gNZLjlO7BDw1Rck+JHXwJHc4ENm2K0OXVJU4dHbV
vvMZjrQM9Kr37Trlgy6aURt3HjlkJsa6ohdRx4lCTPJTOI8+ipxB9S6SxCIO4j8PBXKTajEpZeaR
z8FnWylJSTF2VeX58YmYBNHAlR2BOPiT1lSj2Q2tNMeL1m9k/q3hSJO1np8QGqMO4LGNb3fnPC5D
GI+UvYYjpEJdY87KBgfUp+gJPOJ8U0irN8JPaOjNnj8NLBK/EBeXQ+ECECIaMk6DWiPizjQAlGYA
YV/a2CRtbU6CpTUI5ZAof5z+JrFBdho/QqzOUW7M/qkpZxfwPOyEmw0FjwgBabvaX/tZs4BzG/Oj
YiACOaqZLYBg6tCAM+IgYx7dRY5VxS9rBkbgm3Ytl6/tV58zhzeX3BjsrFI1CSpOSPJQS/6+XLtc
sfvXJfUXxHHQVu4lEAELVWM7/4KgtbfaSzB5P0PrPzJDySwACEbCOebeMp4XNSOLoxCOgXOMqBDc
tQ1XjG9FX2/cV312aQEpd+xeBZSxShoKvr91jEYkB/MkwfxTJNf8umtxMI/h1RcHSQNlOew8d6iY
1vVw3zlTA54aHtB0JAXvAxeRlMPi3glmgaHVaIzSxTgY8oWDxDYEJ515GkO3kRqeodDXrcOhb5xh
2B0LZ3TcIzDWLK2fruwWgf1+UVfmJLxZ0asQlMhApxSEHqp5t9VgEwTzSivFDfcrmLg0APj9jbi+
tDaW3CzQdOF7W+rWp2uObQTdWROUEjscJphdpo2hv9b5XNd6oMuLfSqrL5LPMw2WyKgMD2w2rH7w
jdyfIGWL9FHYYroilmwOIYRCQ0BAPmTaGbuq/wwWHjMNthK9+5JGqdYrPFX5NL6EobCHVLbB75tw
Yt+DTIT0/Wm1UMkBpo7h4N5PoztaiC6QQrc8XCVhwUEWFltSQWWaSMhbUZv8ePEFGHN6DVv5KPLD
TC6fvd9QA4KF2JVOtEhojlL2N/aZhIF6R8Kw5W1azFbNA/C+pqhA2q7PuJO9ru7CAKpdmrRkDEZP
aLEKE1vhfHy94vHkuOMqMVKJlyHx+2K05IULcd5SWMo0XgI1e2SoYzS9JV5cLgSicxal2XNc8vPc
8nxr+x9jG7vlRBRNdInrWLJQ3t6BIO35oT153C/2W7aCPIy09YH0/JfxFV0UG5mXvmAV6xPLc2TX
kKjOwxQuw5K/QWEkdbTGmnz1/GcN5DiZvavOvqStUeibC5T8+iBnLo+8/DNTh5O0I1cxOBLTaBN2
VALrwMi4hwBAxGvPcZvSGb5XNO1xtiTpR5TZ93cakYTGt/96loPbqqmVm89tsIKrB2pCs1UE8+We
5FoRroRCI/n5hQPEdDJ+CVAZBZQlvvcszC+SC5EvJqe57BuPXHw/lgFPCfZgtnaAfCguwLvFgy9/
WMyFw4imLYLoUxYZCpL9Hzt47fNy8VxrSmlQhyl92upz+/trnOR/K4vcahtlzfqd0qho1rHHPtAj
0lvJV4h7KcfNQQz+7BRneXDkiU0HiR1tyOzzOLEHKCAf2xpRHcuxffDF+U5+ojEaCyZeoM8v9Dny
oJ+YFlGsX87df5AS21keSjISgRucwKIQhjldiyvYIWeSogYbC2LlwFJO+Bgp4FfCMkNn8MlHG7Y5
D4tzt3wkClI0bqeqW1hDHnbL/GUTrHqhlcDQgo5kGfZxiqJklnQcNEtwNRYAQvv1Fkq7ys2ClsMu
+i+8I7DSf7TmRRatWlzYsJw+wLEpGnqkfozTUp0a8e/w7SWxFaU8um+69/R6cN+DXb4dalOV0z0Y
hzsA0GTVb1avdbFXubLOWj+YW/ME9DeRcxytQL1FNhgk8tZGz22wDZFr7qiTmwJr1UwVhVL6Uujg
vy0ELXvV4m0HH3eTOsnLXTZZxO7m2W35cCG3xtrFiWE47qfXnxZ1XdUxMy2YtEhuqs95vWcBEU+g
n+uyBZwtFEE0oRja08rryR4wKLgR2bcruqZ6NRjG7eb3gv6CX/e70i+cet+XyEG1yUz70KiRR5z3
tl51fzElMss5FicC5Dc3qw1urjPUwasbQ2m8U7ypXPOEyhQi6IGQV5LJosu9Pf8CmhXhClozps/L
oqcAqc+HTPaBRH2CyY0W2bAK/kKo5/nA0gc+k3Kdaf9qpR1JFsOky4ynVPkp0de0mKbdWLhh1KCK
7H8Z06ge6kMrc4ggWeACukTgnI4oTup9YFwB0p6ntRRe8AnysE4tpjm3AuHTz5HxCMk2OFh2Z6ll
IFa8ZDRrKUdnOQpxIw+ky/4/w3ITuEoIk1513LEyIuGRAgP0Dliuh3nka+mXwsqbJ/0LhaxZQpZd
GkCEZTS8HKtLh8pQRP/0O4JqR4EheNbftZZg2aldraJyN4XvtGpefU5nUdlIgSSJXhXXbT9slaDe
ds/5Qmhlv+A0/gN2LFz1dna1XFChbUVX4G0OWvOlZ+3iE6MGaW0cXHHeMd+yaUQUycqaXj3MaV/c
NooB13CK7k7OTqZcY/YhyP1qS+Gb+8lambAygKHE408FwIWpmaefQm85d0Kk9RhLSqzB+XhZ5rVv
egKsVCY6AhLt1d4hK8mzed0EwNSXekmPSpTsusDCDWhky3JKYDDL+yBH3Yd7tZxjj9oeGG1xyGBy
j8xk2BYP/PPJjLZCVzl534/Q9jyYvqk+h7/dS4XsxQZVElClntadovOMl9BXuVcTMUyS+PBTZKil
j4f7aBZtTMrBG0FHHKfgTHTC2Wx0JxbfBnQ1wDp7OzwPD9edIwf04B9QpT8HlKax7lLz0/TUSMR5
ib5ZvNtwotagWQjBcxq+O0l0eWAj0uGok6kU3z4YZ3muUapoc53dy520441lkTm/LPKA0NLmFnTb
IQTGwGnzk5RCFiCaAuC0+PuNQrr71nx+8uaPBfgGYxOb7xuQvKMFRebYa9yKmwDL0hq+MOe3Gzu5
eKbJ+gKsp5M5si7Ja1FPX5sZBY/S5uVhy9njnkrb0StcklTjQJENqiHkpa0FJKBsOAbIYeJEf1nJ
Ugnu+OgcreDh3eLJ7n3hzOieei5vPLA4/oI7wI8sTUmwYKu+P4nXDZEVIymAN5JdHjaNMpz76j89
AX9og0dQdf7CRC31h0UGycb8w/o4ne30FomeWPNyjaTJUzq0NyeHw34y04cS6OXbWhluU8JkKOP1
+sgoqdNbhTfDaQSTEqgsHR+Tf9o5xeB/zRmVwacOkkmMS7LWb8GKKivjJTN+h8JLj+3zzXo9J0SL
wFI7QaiQn5uGi+/xXqjb/Mh0q7WBcAA/IhmHBU4Qy6LPCyQuHkNl0mtdMuawE3h5GcAJypNSkA09
kxKqZ55PZuJ83tc0yhl7ofHHyaH/ZjK8TxdYAUM3Uz2pX4u1CtOn089lrm3NStSWWV1raLTzKj1B
249G3XAZMLrxLMTGn90/JsnfqCg9CmeT7FHsQFvwybBrMDOGEPtaJg4xITK+ExGPxTjO/nxRaY1K
/H+QqPL0tCi3uEH6cLweRne2dwRh5NFTE4GYXbuCqiq4NK6+4OPqJWlo4N/2aN4xxKzLS4xgZEDM
8qz3Bha40LYzDZD5wbL0a3CZkiFZnrLYKPJkrpv/gr/8OK2GM6dGzVavLylawHQRyu9KXmAqpA2Q
90HjPz+vE6E8CmA0jmyQ3GUjsnsRkcTxcq5MIwbQd+ntSoadC6/N4pu6QuthlIZ7/YaM7SkERr5k
2+tKf7o9E2TPVoWIeqxxDbCl322pL8zcJYEj4Ijm7EIVgYSHPx4gqT4F1foREGo6gIeDchyYpI0Y
npPIZ8dyxuH3CjhreGcKrnFiajf7jGiPFbeTVqnoJOSOAPt2muOxwaC5MNMBeP/Wk4dSEegSB05A
KweQSm57KRepHbErYqw3iaIx387zwH7ueJu9CWonO92Dqupl+nG44IPZrA0VApqHJ3xf9vkdPtXt
S3giUr3YnoVtB0B0Du2bvNsYvAuTTQdTGwAe9/ElXqxQRAL1tloI9qjg4cGIrgkWd1xHszFbWbHv
9OZxCA0rj6GF7v6NUuL5M+cyOLNM9kHMDMckQw8RfxicBPiyGCVo/tVsYTgtSAQoGBax43civbPU
v9AidHt/2oIQka95vWOOO3yQnpjkom/NxkNmgS8L/U2/9vt8+ntPmSO3ie8qLz0a1TIaogQ6eBnO
KUWqKU5hGHx4OEIcyahPiTkWBY0UMqfXUgKLLuIgsLECNZY+8R7yMtXgJ4GIbdm0j/qf8pFJ00ke
LIMu/2mqAqDGfBge9TqrIyFlWDlhm0MncnkaqIvHKwIQWsP65jU0/ZDX4ieMR/IjCxX5cuwjAEim
bwpKFfN7z2ULJoJBo+xb0Y2uz147NlrFFsShG+dwOrn7alLIjPG5VpBATpmYJaqNOH04/iAwjh3B
wJGNioyUEUULjc0AGz86PsYz7Lr+mckkJ+Df1vaq71Ao/XoLUwo+THLvewY6/lnjlt0jrhOeiyR4
13npjlUuc/wAP45TLVMD/N+bh/KV3AwmqJXIi0LuE+wzEmSdY7f4Vj9MpZEbgXdsKVFLtrewKVeA
AKieywN2i+X08WpjrqL/4Cv7cq14772w+ECYh9PhhEVxjSXV344ziN0MT5ZXDIRLbayMYP3QvaDC
1FykA2vzJWvFwXG7VWqGybMultuK5MmxBDAvmtF01K8ugohHvw0p0EBhaozB8ObO1udc1PAhJkLD
S2rKdmW56onr629bKzgGELAADGkT8VHsFIyMhY/C42XxOHoANXY4p/j9GTkpDWCCwDOziWgzBslo
LJdBCBn/LMgS2naRnLdjB+q7wGoGra2ktDmq5w0tSI0jdsQEaqj1xtDiAqEfCJzmNXAog+9SqKy0
ekd+4aJNpFu+Eu6j6YLdRCKN8cnCwVIVZCf/kiwzj3OSbjP9u3mpK2rCvt57kXO4mfVmVloIJc9q
/cdIu8wZNCeUZWVzphClkObrVDAbH9/yovsB6+E5FooXUBvwjfN1EhlhgzAPuR5z8FUkwYEXER9i
OAyd7wLgw6N6i8Hblk8Mj5fj51H5Dkfta70eMZNQqT0BoXUUzTvsTSGwkWyavUovE7TvKZgZ+/8s
LBF4GJVB2zBcXXOAaCZCpA4HTMf2RK1eHDYC0qcm/NsaE94wegKMP1ANbIk83ULmejF70XzxM8k0
JU0QpT9HW5GSHVbO3/QfKTJXJxoHGRCVM5r7UGfjHMeMDRLIm49OvjeEkotwnrMxM3dV6TGqoVLM
s3FCpqsA0yYq7chgbFKwSxs+EX2vZrkih9VfrCa95FFtlkYK6/Vs1xVHSSk90OoQa1DDpK85Ek9m
m/8K12J1N/2P06nNwDSFh7A4Fn5SSlSi8FFBNlfewL0oeU+gkWJrIqCM3u2h28MuPOGBZLroHdTd
gnf6fncPr2Bswy9uhYiuDwLN14QZT5h8KjD8fcgOU2euGTmL364/qSzmaMb7R2QzdQL+RGi/CC8y
SAsEDw02GRsth6VzHfDm9Zf92+Xgsc/N3ldIpBHeEvFsgNgbAVCWOotqMUp96j2I0K2gKMaRII0h
+MVwD8AmRZpz+iwn5dLTJN+LoMN6FDfDX7qXYXYKcMYBwhg2ykkCOwq4wkmI2TtCQMTXoeAgwbTy
E8eR5tQQamcalqLuE1is7km2zq8Oar0P6I3Ag/zDv0QafMBazNSwJufQ0sJE5tnBcW7RMLdYMdo4
P7TY37ZTCxJveHgyrX73l0uoydnesBiXJ0waGKjLNvE5QDswunR3kPhGGXjWKzLp24oHIgAWU9q6
YeM949ejdR/ZztlyqCgxk2rpnXoYPxlkGB/fW+Y8dYe+xkf4oRqIeE8TNmjo+3/SJhWaSpGR0oYv
Syh+796ExU5ygNlnc6GQEiR0iZsseQTRxWyI4lbKE61qgKJJ1jhuIR5MdIpDOVeNiz2G56Wyo9jm
gKUZLoKUAWucUfvJYUq7JDrrRxU9zDR+FfImDiSNaEedWFdYIJaSX+fc0R2Ga9lWkiemICfMLUVq
vA8GbL1sV9FmjsFovQkGt7KIXcVXj5Xe+lTW5/9OzPEAtqtAGMGoJrdhTLsVCts6N2ys7SpWnOT+
c/wGmL62kEyYIl7/zxG532dBtGZjsm6jLGxwnGcrkf7Roev3NCSZViHCdfWqkCm42GR9+6sxEUVg
GoawK4uD+KkHc6LexDflOpFQMsTuGp2UpRQLVIKQxbETnYkx11Z6g74pKPd6N80o5Rk7GCW7PJiG
cdmbduJMPFcfV9RLN1RBhyqeu2fzJaDRWY+34v5SKIVZP45dDkh4clBUZpzauKOYWqbFUJ0JfSiF
PO1B7HBboHGkZK//cJksyDkdN0IA+qFBFUy7ZFg1r7416RRPImhFaIQ+X4ZM8eHceufVxQPL7Gp6
OU+V+XTAtrWhsvt5Ph7mrnfV9UCJSsPO4j0mEge3lgpVWB/F12v7n2gNVGQ6rusqPjWhDwZwHyXs
oRSpgitk5HtP0cbdTxzscZsmEA708VoeetLz5x9tia09MfWxJkyYSzDVu1tdwSJmy80oPk5Nh/rH
J8J5himJFIALBozCnjBvUa1IHzednvoXhXrYPGej6LsDl41RQGnH47HAnHL0oaoUBcKQ1phRWZbu
4D1h2a6ad6MoIfrjuS6GfZc99l9iIzCKaMDu9FA5MPO5XP44JZlCrvJwY8jIUNysv85R7I66r4gE
scIpZijeR7+12hGVqM/XzYIZVICwqRKSFQQa+vvVkoPQUIm0yfjtIf38AQcYs+XRBa6QL0/RHl2O
Uua01lDdGy5Er72G7UqSx+9YEA7lzfmjpUyVW9GUMHQ6/+uJe8vaVv5p0tSPNPG4GdvtQHzcpq3n
lpU+ghuMMA6CP/R4rnAB7RA6ZY4rlw2dFmMJeCQaWBhg/L2MNfZ6hAIsd9ExCqiaeNOFqWXiEiVo
cyrbX307GTCmIH281F+olIBbDk/KrZYKaxlvMKti8EFSMci9DlnDvC3vc5uFLXhJnFWrWgqQebXw
e+X7HQaE0fDIqvcVNNKdT0C1JAwFjMJSSAI279j6wOvkxLgY6UwZedJ9/xSgMiL7X76+8oWjzMB3
ntdmJv+k+2O6MERV2Ri5GJcVxpc9+/zYMP66SnrovSVGfRyYgKdu4acyDvXuZv2qvD74nGEXVd1o
ZbZO0S/36ccrzN2z3QkE/+5SmhGXf4AAZ6ie3q1PcJDa7p4N0xUUVp9pMSj0Vf+zf2/YYMiH5Qqz
bqWwptK8Qu9VM5QqasHOZwCaifN8g5QPKcAfrGf/RaXohaNfIDk5bX54m3mU13OTJj3CFYts8XJG
4EvPtPg7yYZKYZXD+dhJfNay5c7xFtqrv/n4hrUGoWtdIzHXpuPWyyOCrBV6HShYpikD7jaNFFkX
Lkz7PDxx/vPHWKNEwKjklcobeeHLr18UIPQCRovOd5xbgVaYwNq6HQvgkn5MOgUKZKaqadkIskw6
HSKjhx4Mcy+D81P2U/iCQt8phcwI+zV5ornFSJGFZabQdwmz6jAKnsSxuffJi7trPcvB6E3jKou3
xgYHiIgvhaM24+tzH3aK3Nmw/kabKhdWSM8m4ztejgOBM3mNHCcfI8ImcGmNjf/Xpzy2J5LEVceN
4d/62PH2l6QppUyhHDCnMGqq+uaN+x1ekuDCAXtJL+7UbNU9UGyrjd3g+94QaOgL9+v02Bo+VpIA
2fU2RSBnjz/gyBld/F0xE28udB0jSJjszCf8waFRC7lFH5pYjoAEkYACVXdpUD/v62tpFXXHltlB
Y5gcS2UrY/NkTnraCxKpKJFx+DVma0tlJxlRH8pgV0E8o5fnu34OjNbJem0kv1lAY+p0t+cg3b2o
xdeSan/A4SQEosOd2RQg2+J1Tpk1R+DFjdSi7GpXfaFVCVA9wiuBIDM0BGQmfmB8UHvWYnx6oHNU
zBw4qVStu/VgC4+RFz/CKguz49jBzDZEqXwYVmeEtiF6IXVKLeP3dOVyrORqy1BJ41PhInsTOOFz
y2H5Mb2m69tQ7MOcQYjYiWOBCnNIv7aVmN4+kbZHEInhKIOUhHIEdZaLdAgnJj3odzy/ijcNvYvL
mOGqYxYPye/b4W4XYKnV03+Rx0HT3IYAdIYDmlVGB36vN/P68Jq+sBmgdakaFjH0GlcGLDRLpsNS
/lA3Ru3viC4t2vrZmgAKqq8+mH3XfPObX/byivPPBN5Wi+CUxBgMEWTtJEDStWymfUpYv2JxJg+1
PHmknUf9pfRgi4yd/puwBPyqFiRpYcxaLjIig93qnvHecwBLH53vy5SxVK45exRdslPS/UdZqlgX
ac5eJFEHnUvmC9d2w/G49EZwRVaL6vanqHonE00zPmMJcTFc4Fpd1dlW7Ar6exEszawnzw1yqcPR
9aOmMeEPa6m40u+XyqgxB1sftV97lXdO+by8X7MK7uzqAMqTLBfGTqC0JkZkIR5xkJg7g1h0kZPL
14SpzVTmdVzsAyvvN+F9b6EzjONVrc96BXq0c+HPkq6iCYE03UK84aT1ioFNHw3bMjm6edmYjAPY
BmBJjuWj7SbHc/XGQKu7XLsBWSAJbyUgcyBCPtFcfGisNELS9hG6NSJ3+Q8YYFXrJGU4I+lYk/7a
NPD87vj6SRM+W9YWaKOVgmAQR/VwcXzXt23bQHgPDBZhOdARyfKAHrCbsfzkyyyNLFvMO6oN9v1l
kkiImZsuF1wEq4OO6ySdsRdeuyHjmc9cCTR+vo1TN+K8g0DxD7RxyEFoFmLj4q6PclTsxO+Gc1vI
/kVbiqs1NeYlqR8ByzUEbzJK4Qc+aPo6jVmgE7tV27CQaZHGAjf6pVdftNOIldkFSc8p7zGaQ19E
rCroD+hqxeA7Q4wo0Tm+bMMEG5bxsmvEDQinNPRLqaImeb1ZvTiTuOdQJfFyIN9ceWl26TiVkdqj
UJdiezvnSJVrf9SOfoeEqzOKozdd2v9wHgwoyyHOm3SEwndAs4LRKzYX9jdLidYNOScHlO/j58RO
rSHaweovxvqhfItMUh7HfUbSY0E7xIqbWub1rPtXa3RXk6O8Egp6eymf17zegWkqfM5lOE0fQnCj
QPrPZQRSCmSO4AoHFJ2oNZ+48X1JiW/1lyIcBY1ynikld+FECjVGvMS04+/Fcjz35KxhQl3t/DFT
hLCpg7IQhLutdRrD1+wMEmk6+TTcSdzE/1YE7DyEpYyBjY5i7yQQFc3f7uSmaoNbxGdu9gkx4rPN
3pbReZECOlOBexwp/mtatEjWq3SepHdJBcVaLepLRvm/45scdEJftdE14J28ScFL39T3F8Iq9MdP
rae8qJG1vepmOL49Xt6tIUVP5LvD9CPEmy2tvIJYqp3F6B1zJf3FrZQ4fPZPj8PGHmol5EB2SR2M
T5iFSBrTC00Me/70Jb7wdByeSqIRVDxPilrTNM5jl+EnssQjIXHFTYyCLVGvl0khh4PuBy0VSJ9v
s9RvHFxf1xagRVI2vN9tITWUVhzu9J6eBLqf3mLbTd2R+dxXqA8MKPHtG53J5JS3/nOvPL/ntg4T
v43XSY+OEob57zUV+7f3FN0ybqHJPp3SB/CuJ5l9MUJk+bFaNNLqgbal2JpzB4Z61xdJxkdfNaEw
WLbG9KYvAKCXpcBsdbetcZY6uFc9EAaWj7UoiYEsDQ6UlXwctTFYlNng8g4krGK+HBsJKt3qSmWb
qIsELKpT6WpJdq+MZexom/49xW5CKuUiSUe6TqGp3WgsWhChzwVUjRUDC5hEiGDgGOImEGmphH67
9jlY+nUyn63tOXvLVJbn5ESvcJX6ye1vVaGNtpkK/1vv+WMU3CfYt4CaZ4vpdyI6kJwuKK0Mofwp
S21UZ07L/yfKbjIG3Z0zQn8QS9xNhesPwtqvN6HYjjdbyk+c+gKYhkBcBiTG1zdC6cVH/vRQ4nw6
/vN7FX6qaPigHTEkRYDfBO3z+pZPQRlt816JlsorP+Dn7GilT8AS9N5LzTNo8aNRKHkc3UvvtsIN
SFiWgSzu9znL4GjS4iwLvg5eplNH5wQ02nc4h49N474INmtO6+k9KnNnH70GjP98QAlc5DRLYDFc
bclPW8UTav41dTTE/KyD/MxmcZ4yNArDEFvar7EdEQ1j8ctmQDem1AY2FBdEmpxb76HPzrk9E8uP
vCTwTR+tt+XK7yru9ohR2EBWCK0IcEIz/aRkvQN/xrMh1IIT+lbnXG6U5Mcd6VSsw2TMTO49267y
BLTc6fkNFixQrWhBSjsr0fLxYQU6w0pbpqcHHJHiujaYFH5A8We3wNBePKOneX20isw3PQ0OnsVR
dH5+JXl36Mo/DzUGmsimr7xb3GyQ6KsNedJrFc09jPLVhH1/eWs8jE+z+7ahcuiuvG7rawPThGwx
QK9TnP+GQ0jaE+W6RFrJKuZaigrwIU7JA0qvIGsY5J+iry5bM7owJZj82F+ZF5I+L4DbR1cHTRv4
JmonAKtOxOQzMM5qtbPwQ7vDCKXMMSP/uj5l59CbEcicmypii4hdKIBW7GhSJoxdDQINALRp9nxf
2hUx6l0QtAkfp0UzGAul0uvDCd2hN2vbbF3NtZ3Plbhg8YIaiofcPI+tS3v8WmYVaWMouGb2Ucby
ohIzaoDM5pgC9JIHRy7UfpKmaXO3FVtzsDAEWQYCQG+PhFXqwdWCxAKo9msVZuUQnIue8lkq3Ss/
24UYaNoaHpjjg2nZk+1MOmvbxMahrKF16c4T1o8bh9vIzWIpsYZtdtih0YahGUisYfG6y2xGCxYp
Lj1tFJ0XqqHqEIV6VIwJWL2+j1zRMjC+4fCwEJnXxkEe0dfQv+SxqAl47HkuGyQVP8piZTAFTxoj
HtXJF9vrc5oJdygl+oTX84MaRpo+aLswZWGXUT+09PdKQQzzpSWh0lzVnr0wngBVUUloD/npmOnZ
Q7y99vYe+3ImTuzGvO6KXE+YN0rSRZYtCCFA9DOVXlIb0hpjuy7vRk5hsQrgVbw5ROFmMuD8SeEA
40q91k0DPLKpvEnRwiWBf2tpv8+UzabYVBPzBbyYIJr+zay1GZFT6IUKG4Pqs3OAiLLsI1t0HI30
RK0n29F1d4FUHkC6ANjNL6WACKtYTGgPL3lJwW1J/HkiemP13MpZxSEUbtXi7l8Fg05UHAPf1nw6
SL0CHfbdSTOxvmTdt3L6mou2qidV9+wPdN7K3pTym00BWhq1JQi0/fKYZ7di3vJvAVHHTVqCVBVn
C68TtNFW+xobLB2lHn44Ltensia9T96m1E/VUKsWuEAX3b0sqD9uUnssQP6szrc0t731h4kEyEEc
dYzoSJ6/FRcn+wYqWQmMY+OLZ+v3k1YmZmZ0pSd9znYwWQdXcafKFjNDPVNgWjwEnSILQNtPxwYU
RwOSzBw+9n2S9X+rF0azu1d7n3/v7vn4LSCsu+opgrmf2766VqbWREQI+b8qcqDeZUq9yCc20Xoy
92BshXVEdke9jiZ3cTQtY1Q1A5Z4m9dGS83SHWsCMD1fxpb48Opfqrh30vfmc4W/XPJZEJ54/mZo
75MyltKXtQEXxDAj2W0p4SYetruOCZG4uFqBNrbhb4WhW5KuKGKKVpHRYdeWrtpZ2EAesDPb0XN7
Bu4tPhDToqA0+Vq1LCRNOW8bUzG3c0UT3pgXYHxzuHWhXCUM50aAAfEFKrH2eV6hlIdG16O7DEuF
9IF3/O0P1T4UStysKk0HhwCAURjpll+F6AA3xAp9QICSgGe7kyekTBTjqguGVpVYbkDWfWiIvl22
cRHV+LQzC9CAcA0kkpgHeVUEJnf7JU4NlSHdOKqr9DIK+Ah0T+kU2cxwjo41tZUbpRJxmsZ4YXHA
bTJXdsJRo+wB6K+7yhYVaajJnaaLsAmoYuLxZwxqL10ynY3jh19osUr1d6/e6RWzndbQ2n09orK9
nSjRzIY8l4K7e8UNIDwjd4ro2pmkvkijPsEkK7bBzhVXeRiyZdqV3uKwLq2Phbs7BF1zEBWht0Kp
2ylC4487Zcz9y+zCOVwxIKK/DK11R46O2jux+Ug5OWJozIEimDZgEhVviP0wyHqMHL7rXU2ewJQx
YW5Rpa4tH0Z8yGhRjdT7s2ICHMlA2W+TLjkOwjCgG+YvsqtStBdYwnz35ZgjbFCSu61W0bPxewjh
u/hTPDn5gDzjFaiWyvJGthVJaDK4DUs7XF+tGDn6PWDDUjBKifgtZEbyX0cAXjHFulcnCzq0m+80
NpSIZtZYUTGcsKhd6OcEDQUCqwdv5vAqAGbbF7i3nP+xnAugm3tWyjBidXgIuc4XglxVwIg7pR4y
71TmfC7Zu0wHhmL99w6UdKkwV4Tl2agYNRxHlY2ZxPCm3yOFIE6fl8g7PEBhRFkRgPn705h5d7cA
bd8bClhCEH9HJQNuBwwohYObUyYdais1SpaelZaW7GnHxW0wr3buGV+C8Eu5JfDazvcRYP1/t+im
mRtByhUIXzj3ES/ElMmkbF+qkt+QS3SY8tuRZem9d6U5vn8mCR8Jau0MQCOXXhZJNhLvWEGRcY5C
VAYKo1JU1TSmGXsKbSBkxaVsF7RSdQOpjNURMkbC2ojWqiMK47UFTdBYDBw7+8+SYhDVy9jf89Ch
Jr983s37TkqqCM0eWoTR12+E83865DJWPs4hlOPgPihBrKPFGhL0USmPFt1yrZ0hXI2Jo//gnUX+
hkMOOapH/fdOm2qnbySzgorV8hFoAjQUYmGw7KbPxDuGDOqMgKYbUMoQkvBiyJ+kCAMDSapD0c1S
BtkGu/JdxWfGwX4kY0Szyv8NG2cex6JxtqzjMa3Xux4a0ZISLylpYwf8o52PSo8XddZt3gwxgcko
1YoPrf+zlsgQ5nT+moqpyn3KUGylQyVpuaDrizRLmcvm4975bXK2akxXqWbq2cfxDf97nhLRRxLb
BnavdZkedFHoQxAdTYFsdMDnEQfu2ECMylvzyVP7dqU5ScUKh7t8qwG+/P42q/bkFNvVmMtPcndd
GXJRipXGPxt/Hyw5HAWfzWlH+ThJP4BI17bGQ6eB+7s1ZiWNSHcCJO03en2tOsn1dp7symoPPnyp
RL6GEVSVly++Yw9yY0ybcda9m3/Yw5xVd7lll+3GsnoUO2UqBUFjPkNP/Bve9QGM9i4RQMb2FpbT
bluVbF25Y9kbklqf8auXp7xEaNR3d4O7Tc/9+i7MSwfJprck11Ynb6tfZJrUaZF4QHX+nASz7YO2
B+M75V35y1+VU6kjm4IvzJ9pY8e6NWv34M9ufagOQtbOnNuBa/1A27rocc6FyMr2GIbhjaeMcAIa
ZIOhHkvF7TFwxAsU1AeB9OOU3L7/PzpOM+0BUheQnkC0ta+tQPTK1g68rRKNFsEMc1QkTAqhE2MY
u7hdwDk9QvpOPlIQh0YHtXKEphDRZYd4NYP02AMIL31BSSD8qf/07+yFZF42S173iQOEe13ZMLDh
cx6iLlGlfvWmf//jtIZxXMHh9ABEejVcFvHU9bEfyWgsCz8kQGO9NCmYGcm0y88wWmid8tHPYenJ
gN9n1Voc8PIKzOiQlk8Ev9n4+QZcB+6qN6Ztgu+AkWzJPzCpiZOpCfiPZPLeXHAp+tiVLLa7HIaM
jY064wDXS2iEqaQvBA+8ymu3GLf80yc0FYNqsHt/RnvbjGCumRP/D4KTAAoa8Yv55UvzxrAXvdYf
53BaCVxB8+TMg3n3w00ijxx/nADMuTqIj0BMOI1jrVRfy82v1Cwu3A+ZXxLhlqvdPpDqq6sq/uhE
PVNZOtJoq6QDTAxqlPdexa+0bc0sRzRCd6CJGXaGtasurwiRsflARlzS75MxsjLd8x0d1S2uPDoy
OB+t3J/lbAPB+7+IdIEcrUvty7hYLkTUrNVQjwYNxO+ePvarOwye0UORrNMm4nwWpAbWAl8VB83H
rlrt2AuhNgCjeKFohuVYD9xnZU1e06U1meFF3O6GRmQ9B65tcrNtfmaLa9jZ0unywepjC3YEnIVC
2wszlD3/TL419QvbfjIuj5iTlz6BLEDE3rofem2AFgW7iHJ3FPl4o9qY1CdCeLROh6RtZpKbp9t/
ptNWewLGm/ao6wDrbHTlOozJWNCs4BdSEs1mU4x2Ms8tG7v+IitDxtC5O1FjL2HcOh4SUp1+KN3R
/i57Rs6m2PxWIsy8PjvxwCFM1CuolostPDiNL6sEXqDXhP4SXIq1JSjpO2JgeH+L04Tc2591CzQ5
soO+00JQvE7r6Vzrrs4jHKBQgAaFv1wTAvyR+gd/6U9KrEpYSfyNF8BW8qFsvQLCfAOM8h69quyd
2LGQjnr1PRXMuLAiJpTOVpNEQ1/v6z88Lyt0wNwWpo0G4kTcVSE152h5IIHgtzglqp4YtcD/GRKl
hJFuSFO9laxpGBz8YdWXk4u6vRD1MVn3tML5plO9tg1ekGzNPwJZek50D5nddW9Qvig87NNXsyUy
9zvn0lcmDNpx4sI6x6HMrosnMuJIpe4nvYoQxPmJfU9E3wD+LhFZssTFi4B2sGINvQa+h/BjbA9k
b5M2G/LKEugzh67LRin3FposYii5WYYA8knBkcUzZznHIH/011WPlU5Tut3fwVWYDu8NL1sBsaWG
TDyq7BeJLipQPmFTBB74GGEwja55nVYC3WLw296g0HSyGgxqeksCXutvNFj6tcn+NXIJNNOmPhJR
jIcoS9+ioFAjzEBnMaKUq8XN/DWD168WzeA1tfe2qI/apfjRlcBPRUCvHZ8cxMI1i/6f7Ly1zejb
E4KqHq0FNHniUPqI8Ttrs+uwXMFcZHxWWCjD10TcNg+psWaQHmJlP9Xolwv4Up3TnPFVWfOcLuQf
38xKDl5gGZ5pE3XeiRzJgeNx1APxcPFNOHqXXM2/5UUt1VnQPJjxoNV8gQ0LZaNKzD8ILQuIPjm2
xANaa+J+QAiBaRARz/g3HhwoIQ2vB5DcIt91cc1VaKDaIksMe2tqPWqjeIW17CDS7PrtQUmuuMXa
Ti9i7wST33pNu4ceczO2a0w1L52S3fU9Go/HjB9yq9fNvaOicKq0FoHE4mi5xdJ872deVCyTbry+
iQX4eTmtgdKY6UM7HUdcFbuzKJW8JXa7+51cym6gaemJ46C18XMFzrUgdmZJ5R6Ii1nYwu5IaR7J
Gcyj3laBAyopLcfpxEuovk7K8FaA7uPcjpF202/D0z70BKypeepIoeBRMiCF8fNyHZEj1WCnz/1o
L3qd404Nm6OZQEq0FNZ98wel8PaVzeBRyG5ZZdtTtm6+GIGofxKQXN6/NbY7KMxdNJ7x281K2xgZ
buSdy0wwlbVqXLvH+Fx3j5XcWpzlbYw8EG5Yp17rBB6T/x68KiccUREuvrRUKt0rLXB8y+FX/1cA
PUv3ec6NXseYIcnTa41mhDlIH0ouWOkmJJOUGiww/z6JRi0xToDp+zXwYul3QaMTbwSkQlWMMBX4
51I7y9K/jfNSlsXMfOM4PkHBT2OnC5dY6tba1+kqKQVCawfgMpTqTLLHNk5vUSY2PUxtTW2mRmyA
bglLFZlaezLZANX82nzkgTigmPM41+VicbI83kr/afIgWVogunvhhnqIlVAeeBt99PIapEMOafDg
WPct7S0aDCpJSBVpSMLsQMk+vEheHjJlbf2O9nuKVzNtIsgKckAUJuwERnTl9UsqW/o+cAgeLmD4
9eBkqyQmBTVAwXOJml7gql29WIM3o4L8uKrwT/MhSLIvXXt8Cxc498z6N7dmAH2S+7kbGSU/IhOv
jAxIBSRIc09h96hpTanAABf56xTwyK6eDa6hKST4ofx+8P/2gIDNLJXOc/XSj2rFMwIserv5256g
Xh0gLPF03AAhy6UGByMhlTm2xC3kNwUUZQlHavt1DLd+xEeIlTU/EHppp9iQKEhGhYyX1yqB1CQt
JzyPQrzeHsD0zBoBABTs/ApJUwkee07HU8TigsDqiIdKT/7yOJjAOAEV0PznPBN3kE7FGs2xib7u
LfuTv0IVXYhSbFJyp3TS1KfU9JiK1umTSDDjkjBLsBEaHqoo+3r5CJBDdMGtLgSM+qhe0quXQp7X
THK7i0kdZsxWYIgjK+OeYijw9NGB+jHOywvKgsaJ/JufOW9KBtVs/NHIjtuTGDFhRpfu6bdyJ/M0
mYztBCZEexQZeErTdT/AmAFJDOaN76FgcReCudTr50ud1EXE/p+z0suRZJgPySy2JUsaNO1htGMQ
DyNLGSTlm2ksC1kr0LbW/Zc73J9Umdb/3TAwUiLq3CHQnyOlNQnZByjz0xLlkBdwH2xSWmwR92T4
Fwkutn9pbPfImQ0KNM7EI6V+QcqqRrzBAHIQQNdMq6bQFGB5jtjqkdFDeRNJDYV1rzHBmG6mLk0A
FNtz3phKxFxLoN9kfxQ2Kb0BVd+AmOSxcfFPuYWOJGisrr+TbEr2HikFdC/mNEvrT2fPJmFQ3f0d
6iK0nH179c6HMAJ54XGsLn8PDWUgE9O8a4+sycBGi065EG+VVVSlPtxm6FW8tS8/tI8lrq/Cnuo3
YHtYje3asDbA7U8kkJTmSG57pZBCJTOoYQvkl6LBxCV5KbIatDW0nyliUzyS3Yut/r0l3nGkS/IL
iHAwyjleG+oGu4dfMm7pWFnFuxeeJL2rekYRL92FZzaNeCcAcJStEk/1CHFIzutMOJdgVJeTIXNO
YlYWVyNCnK+gPTTrzhEH1qFJAaaZ4BZ3/AQy9wUW94t/3FnvWiH08ARA6nN7hmUhpgJGYBRvFfiA
Oa1uxlWvvXx9Cm1TGfAwg3+RrESRlE/uCDXgeK+P84PgaLFIaFidzSxreDufqTcyVrSTgR+Y4Tlq
x7KdLz30Lsm9qPyN9VkglE5wOCKKafSCAvTplkGm9nmoKoWT06s3Y7nlRpefXNUggOCLyOjW0Q13
t0X1wJrklxphOasBZn0PEA14pmE4GbhymQIZ6YfTCc+pbTdsayepU51Y+HP2IbNqVvD/vPUEywgW
ZaH4Ks2fu8WFNB78EybJemXPdeVGyjHZoMy44vIkLl3n1b+Fw09JfYxubYyyUTxZfZLc6Qkyn3LY
AnkjOiPQndxiZnaWggRvWnwpVJH/hXQJ/O4QCDIMm+qPgJgBrVHmxInv2OoxSIN0S7ZDpMnuyMJT
YlIQJGHHTi59dRkWmpMWoAgXqd+Gfkj9Wv3ek383zKY1UkdYy7Fg+koLI7tcl3Yt8MIuDnK+09J+
flo3tKiFVFZIKmEkhA9tubkhYZ2dS4ZVZbXeZ/sMaqDyb2v9lXTZYzIHNJasquACx1LYO3KUX86C
VQCNsxbT9Pu8RV8me/IZrVmUEP9Fs8SYqcraQ8GYA/DSJZ3cK7AaYoOyLBJ7mpms/BrRboHZ0/5y
tNq11+bZ2MaZk1THpHGq+OblE1hRCpdNbJPlTLaJP5+V+xk8cSCUsJu6lCQZGe+pkaubuRSo/vK+
S4uT6Pm5wZaV0s4Ix1GmTrI2uMwnpZVZo59NdYAF0GENo+WB278rf+E75yzYdkoCorszTkGYVH2l
9MX1bsws1/j9KTR1SAddjvLB13cTJMTILMqFdKZs4RmJRrS+1l+/kJp+MntyTWVcFDJQOy78OngC
OQcl7L/bcNlfY5qkhkUl0KUnqHqet+l+nvs+Ef4YMI/RyqByoNfytZJUFI1c8UgWyliV4c77lV4m
25ZNmpwrpETRQSywRDkWDSFB+UMUma91PsinVN5wDk+CxnsYJ1NY9oLwCh9Imzox3r8jLgRPZ7WI
cyntyOpn5w/ryoe5lmUKWQBRL0ggCbal3keU5sbLyaj6fsXaq1/OiCaMfpWn2jDvFw7xX/stZuJl
T92rJjgWgrYkyaCQi9kyZQZH2eoO8pUYi6JG4LNMsU4Z2MfriV4MnfTaxSvs5oZr8np5ZpxYDMaa
s0iP4UEE8cIVTZm/IU5KRB0cp7BTgT6x9NOEtQfkBawvHR5mdikOrit1QB0WbHQFo4vD1PtT0ctD
/aM7S1clWhrc30NAmfapeB3Ufg/Q+UkRZzMlDJajYshQaXvFzimxhCc5upowyQX+W65JgUPwiMoH
4r6YjvqG621UhdblNM6lRgxGnOXBPPOk63gl1QOCMhiqChYOO0zoYgjwyGt7AwzXcIBSxs8NM3ww
9q+Cjl/8PtR5pGjBeTtMSUBULjbX7zmnyQ5ks/2ZrB4FhftS5tvQzcn6/WlEgF++OaIGY/M7YRGu
cEBCr12XjS4PKiG1voXnBvtRGj1UrCX3GnsEpI24Y38/BhfK2GDyvhrCqSrzsbCjw3LDGK0ybmGy
GjAx7d48sd5PxYugvTTZ6c7aAaAhs+qD8UVgcCcmo/gyw/ccXA3jgFlfXXxGZEClQVpZ/pxArG6K
svHF3E9OpgPuHwxgnA9n9hFgwH9pGJap1FQDXBVbEAU41PzgRZFum2IND9jUgwTE+eGCw+b8oRsR
ZSVTUG27/BuH488wXLtvLsoJhd7W/hq5mBghGKS5Int1nULDFNHFn3ZnBzn2+pfWeS7u22i3z1IK
a7qAuvYSMzFdVO8bPjlMzJavYnNO8CF/uIDUeAL8GSYNssgqmhZ4k6fQnqgmn0uxtBF6eCZ9EzJD
yN6XWP/rK9LgolCgARR6IypgXiY1LgCtMRlPkJAg0zESKoiafcbsEbddrBFZFkplfqwt8CVmiea7
ZSS0dNfe8jiL5KuP2MOiOv1ElkedYZhSCD+ny36nqViuZ888AHaXDqpEWhuFiNw8qGKcMGbV8LkO
81l8utujb3MADxcIAVTtNys78KgDwGm/jSyECTRVpBiFYcGvdwM9PbhI5YE4hBr1HdGpGb8+0U0P
KcpdQoTFl4CZ2nqFZ87robB+3hcCMf/id1FMOH+5+SbHAsM6ESWDiieTlO70fHJ4yaE/ZE3Bl58G
eYHF6mNisiLH8sMcOxZvE1d+vyE3UoqyBHhmqN9wkYAG8gYro94Zc53FIIiC9i44dD8xC1WaCYvP
cFXqfTywIKtEwyhPOEWgNY3SOKY7tuVm5eCFc2DqEYxVlLB+0QdFbhsawBn0zk9y+i1VB3xRAE4F
Cf6coEhSe3Vz4Q3vDOKXH22hxjAish9QQ7rgKB/TijLI2jp1ks/FTJD3lYFJPcEkrrRwaE90Fy+j
hXMq7vbmW+pUOUy2WZWg8npQ32IkXTG2G1T/Ol0mVxk3ID+9y9sJLQso09cZF2d7dW6xAG97VonR
znWB3n7UdaSy06qfBXLSVZO6ZrmEyTCR8B0cnzGOsV22bjYijf3sjt1JGp//23Xw9CXRI0sZEgIF
dSXfN55FjK1tDU6AO5VlnYmrjb9LotIRmYtotdZVDHIIa/QohqluTa80RcmEt7v1eAr6bbH8Qng6
NSA+IDu0GEY8etI/M6Ufe988pD59iQlZg3UuiG+1h9vuYww7Uka6D8D778nd6FgC6x5bBc7N49td
HNv4s4Qqn/plDApcqY6qnj1708UScdalO4BjZrKAWfj6NH8LyVaYzjKuZmlCi8enrI2bEfH/fWqY
g45xs4ieWSmxjrxMh2VdhSVYDh8GW6lREyF52O73Zk0PMKuwkVl8fBEBlbsu3fQUb8eO2Z4VKhOP
BbSG6XJNlvZ/56ghilpA9Pb5QjsZ2ZMW3Ix37LEnCNOuqb1FMx/eTNyKVHT/FgBN5hHA4ws8GBZm
Z5iubDqx9sXmqXfRyd8PZP9X9mMi1tUsLOE/UXc2JMEr5ioWCbp+kCBQmzJfnAjVSx1eWzzKn3vd
QKLw5NNOo3AflrAjwFYD5JjQkY4H/jWQkQnMw5jUeAqhpDUTePphCpARb3PwA4YRHkBF4q9CXPAV
Eqz4JIdZT32kld9DaZpqEGpo5yPA51aoiiWAeohAwiaYCoz0o8ReTx/0iusFlFvYPxnQBxTp3lfs
/eYGUJVCVtvFKTMWaTfJsdNKgUkjXVzKkPu4QuYtdo09nZdGDK7LcYwPG/sO1sieMJO78k6ZcA2Q
H5r79AySW1ggs/cWBe9M3moqUeqCfRruMZNK0tHqGi3jNwYTfVzLHzFuBNErofpdG3o/bmIFOcjJ
kLgbSW5d3ATfTF0bjpAV3Es8J7nXxUhqa1FBQBoWRou7LZsGrm8m6yILcrrTWSfzi05Npvr9Fq+A
bqwnvLfJDTi3LkTYI5c9Fo2DOKajKcqsUEJA6PDmnC24FWBBerSA/1wzHMzln9TtbWdXmbu/pUcR
u7RIGLMc2eO2UK12gf6Yu79hH6Zogcd60Td/de2yWoDtwXW7kMrdtlenBWRXq8FV5ICzaXLbyb4I
ah0w/QAeD3ZgdvuBjMwThH5COG5UChPiJ2bnjH/dMQhpjxbANhNKrHW6shm7wLvGlLZVu1kZzCNV
QZ30EiLma+dufMN6oeq2WNsYUywgkCR8AhhF7/5O2x3LOR2Aq+lNEWMx8f6kQbTNV6pvxZGzsCc3
eheBtBDHwF3M+ecSPmcLeu8Y3brDrj5bMhY6+pCtDdpt1nsnRtXda9nbouVUMsbO5HQf6iC4jqLH
mhbb4v+YqSgxNbG4RbhVx1Qvuq8vxgx4J3gYEDFScdM3lDS56Sp+G88gWTm33dUghzjodqvxvsNr
vMIljKkBGfkbOJl/6R+Y9yDlZ63AV7pK2lpi2TB3z1gPPrubM6b+bKY2v6mWaNE+yZH/sOuAMCFL
zmDkfrP92Vx4AO/g7Hps44wnyemeqDeWYARfAqVZ1umd9LXTQhfau2Lpo75GpvKwrsnUXOFeNuoJ
WFbcYSvqygvznQ8l1X9iCGUPTs/YNWHlRgUFg5Rf0VlFjXGeClCyMF1PKg6nBJe8UzcLYx3sojau
N7NQbD73p3og7Niva1BtxGq4LJ3mo9gkD6NZYhe2HddhWq2tv1UPTmVyw9qiLOXHKLNbyEYTYCgO
41QvoBELNIDPX5vU2SD/8Q/8H+YEvMTmarqFKAge9lNkPflyFjIrU07jxnX+IksyvGdflKZvDxhi
pc4wv+oc405/T1JAnkjMTHtDT93DaFXcPnMKEEkO9qEb55R85TeV4TQGgLInethoUn/B7WQ9gD9s
vtATlRMpTGWQFB89co4damt0jVqHc/lON+ZkCEbLftifRY2zXBmlU4Ri+2JMj7oWMntns3ZBkc2M
+ftyGjNCc0IA4KnPkl03UKOOnawWZ8cXaSF5mfaGKl9C4Q0WBWUDDGTjNsTZ96o3vC81j0ZZ528x
gQQwPF0ye8Z54XfU2bBH7od790u6HzvAyNqVIPEaU+T67EdrV1gheCNdvdyKk6e/B/RrcXtUqgRw
gNIuOBZUKfxnTIYDDeSxMhG5NJvEj32s4gG+zRu7aWO8jhbroiCWdSHK8Fm1m/NeVTzOGNB18d12
NoiPkePNh136CrISsK9zaokAG6SmamG+yA/6TYdaYHqk9mSMIvbLwkUJrjcvccCwLijAuxeUBgFb
PlUDUTM8FvDVLkBlnW1lyCy51gNXptKOr2/8+rDOq50UbPXtwBb6qlKOyBa5RV9Ld5gzJ3pfuDxd
x0+K0cARGB3Al8s0T2ZtdGXGgDVkYlJftpHhvvIdK0rOtCbLS3ztgVymCDEPC3iznEU7o+BHkluu
p1Ez2rkrwGt/cwj+Cyb8n3EV7DcrzzOIOQ9C8vfRGOZbT3B3FNl2X39WPplhMpduuFiAKRtOjGUw
wRj/B2kJfSMGVNrtVeGndfJ+sI/ulzgkacBBdzQdkDPPsSPzuNdwxid/YGSbVQ4Prq5u2BhiFa4y
8iYaNNWpkGMSq5/3gQWctuvLkmmZp5KGvUrk9FhU2ta3UlxahqFCbY0r1hDPT+SzkDhQnneArBsx
Uu6cucfp7Yv8enRh9gXGDTpLfl/oJIvSYq62q52HhGGdm0MxL8RqTh8wx/5gU4KU1rj/bfIHl95Q
XA5fkhmZenB7p91v4dTMp76mvRSj3rbwmApCOZpatZCxjhNF8WKezU+ka2uEcykezwdm9J/3jkef
knRxWqrJ3dqZvk4wxWpj5NbI3e6JO+A4B6s1hKRQ8HDoUL2svH/ZYspMs5+ua5sjPUNzVyATGn5o
kovR9n/D3UeoEMDkVMpOneJbpAeKuyzO5VrccqquJcvpoJ2wtgx/Znhz746/0hLJLx2zwVgUaN6M
EX5vPJ7psCrS7Kltyjzs0qByakJWHhyWJ2kMY0adKZY3JUMbU12fi1bQTSbWofmmd2O99KW3j93b
qYH/QS9v1ppZfwfE43HmCGOcbTCkj92OWFwwtTI4y4ZraoAKdi6uL62YJ5aC7jxcdit4rqSGHd9Z
x93S3CCFpk13noIxBisqb258pItBppnUDMRJfLl1h/YftTSGpYfv7Pz6LZ1liIslFXrTO/aB1j2I
9jldJL9A7u8DabTuszhEBvyKMzojkSuUSUehGLU8LZ6DtWHgSIvPUwSZGrHRAOjs4oL0uJhKGppM
TpfvEGLKzzQbIrCGT/pD2VzQ6LDi92fbahgzfFdzEcZ0qpXiUfP63mON7WkuVL5nJKxVDBDZo+tY
drrDnoLBaGby055ppZh8q/KCsiEZniq0eJOZNKilQXPL6sPCZWuo81h++rgWD63JLlLpCGfdZSvD
syLT4+rkHbNUVV1nGF8Xnthna1CP7fd6izl38F2gka6LwAIltblLfHfQIbliSzEkTzRa+xCfoYwM
AWbZfkYRLUKlzyDlm6seLEXx0oWKbWfxXcnsVdWZ4K+/kEPhlBn0PF4cP3GaNaBzbtP4xM5lYOkE
GX3SNv2kJFrU/l5qby6HAbXkmtmiqbKILngKY+4a/eYhNLXPyaQWsHQH0zl3hEFUtUVaag2f/z/P
Ya6WWn4G8SwTMdhwZl9wewFpgCUXOA58vJRePUZVaky/hgnjV5RFugLPz+1B28GeRNtILc/TPKTP
dVkT/y7069Evmbnc/kwJz9CWD/4fx5ObjzZ9ocBWay4yVmPS47O48/K+bJhX9BCGwFGDpzbmuCwB
5JdX7ETUCPat+LVX13HFF34NsHc7zIub3ZPXFpDUWhGDfDOIQ7xRxAq6TLhfe0p5dz/jlIF6PkSq
wUZqWAl1vhXp2VY3OsXOxhtHlKyXymrwRtw+wZ6cOXGaID3g7MW+Fh/5O880umf1w5gOYVpwUDAB
oW8zbvUvpmDznDgDp7SuIQb0xeSsMljFMQpFsM2UPaNPfQFWgq4VPoZDbD5NLvG7atar0+DfgS/f
bm5Y2Sme2bVve15R9ho5OSvtlN12wTkgILFkoi+6s1HNu1k/yXPdKNu6QFyDrEO5lbS3oMG355Pu
gL+Esqkkzogqz/4N8jhmDpzE0jBwRzol/79hf2RbTOsWs9acj8ImuywLof/2yCIF53fO1O2N9uXh
84jqGJ+Y6lWy4e6qQykeq3eexKPJRNTR7aFbNoI+U73HHo7P2tzU00/VTRZPsmX/c3y0KChJ3pLM
YE213QwmkdKR4kyu/FI7h/W7Ojcfl9UGyMP1Cugv41mshoYioYX0szbaJSv5OpAMEQbscZor2Lr1
GyTF1EJR4JqnFL23VcPT62GlRRxoV+/UXh0b7BYnsIpF1yLLEGvMmq8LfKKgZNiNrkuwJeZz1uPQ
wOXz9XlCdvTmw493vfuv53g6USenVIH/eye1mfCLm7lkD2GMVjPRRcwoft18GyoXlAdv9jEXXom0
yGzS5SzzJr4tburBC0V7JAoZrpbFWZoL2BNDNEkJ4i3JHunGLJa/3TXJJ0gbqtyMoDlsd0+Qe5J4
/aIzcqt+jNwpAfpjWpZsE5RjpkgxTRtZun/k51JRRf6iO+jxi+FFSlqgXY+KwweZ9zNJeSE2jSF1
54J8C2ryEl1P9K0QlNtM+M+C5aks4RAkRcv04J9dcKxAjxFd3VdHM4veglmYs1RnyOT4vQz38Hzv
lq8XpSxDV8EXPo/kqkzcdvbC3kh4iQnU3bYBOFzwBsKacvhmRGKg1HBxTlMPdOqVuyTDTLVDiIjZ
Gz6U7oLgBx7PCcyg6vZFUBRAaKNQCQGViVaNrozS0nrf/KNO5m0O/Ulc4n5UZBV+2jErVgnuUIeD
zPPlovhXANJ8NsP/x2I+EV6YT3llJ6TUV+pD6oUh/eJ9VgTEvFJ+kjiKQwtaATZWv2sGf0+lM6Dx
0WbDueVxB+jrdXyIBuh1ypMqjRMr50Z+PTjeCkIq920D48l98m2QkeQSIN/3WNNcIEU3c2HsQ12n
YWSIme05O6SGQVc6xg/6KLsBRzOi8iF62/yqUXTH72nYtWVj7eZHDids7FYubfMNrwM284DAjQ5r
vohhgxZFYExmLQmmimX0Vp6GsBCumJXPuCIpKx5wpLQ8mQ9Y4dhHyTSdoCV2A1hpS1Rw1nCt7wVO
4o5+h7BvDrzVD4mjxgHQmWAuvlPGf5IZi3jDyUUcODI0v5ssNifsDUHBFSSaadi2V2UlecnTVITO
3equ9SV7/axTDzvLwoD0oZvbk2QvPkxQ5WqbEActvNw7+MT9Pi4F4Reralz/8cH+1nfaC0tFtITy
PxX0FtN7c9lhnyul1T6WhbUgdVB1x1Ohlm+6B45PzeYndPm1j1sgT+Ific5HfH67a09/A0iNKvpp
wSzBxPEGR5PDNRiigq3fPWf1m+j6SDllvV8zgmV9wsdqxWEO1VfYWzxW24299PDNvqyQ6QL4spD0
k473wbuqm9L1Ox00Jy5cLzsaPuL3a3obtj6k6s37uTX9WAgBRYoQ5GIRSpwkVPikPfIiRvE/TvGP
rCWl2Kfau+X10yiqOZzL9O4G9AdY4gP7fFEVIqHt/shhTRZPKHI62YFe8U03Oky1JknsAWvIY0w0
r7IBgpCLDsV5Kw2T28f9oi9l8vXBgfPzdj/klHoLo58m34DS8zootowirz5WlomFATfDjCExaKzn
w3AQlo9PVor49AdFprFySGJOa8NxqTCoJLr3WdC5dRJapkn2z0X9LJUpeSCIM4zRx1e2Hqfyc1Pq
/Uam+aL96yoG4mw99E0ehLN3oosVrrcp0+ChLFGG3Q9qxU4+v0UespZpSkvEeSMOXP1rscmRGWdw
H5CpMUU5egRha++SR279G1UocsIMGog6srIVs/9+oBBm99tkQV+owwWpFMF6Hn5nglEzV6EIUKaD
gIfsF/ssqayW/auO9UOD+n4B9v4PP5KtqR7TrfzzqlUfPoev8RNOg1bMXE04cntnlu/yDv2EKW0j
P8opW4FXKXGnq99EfCyVpnHkd+b4oLjkbiyEAa0OO5/s30V0FofAVvNmosiTTTLZ5dNh7rYRCnjF
CLTj1aMkYNi1sxQ3hrugY6+wShOzrRG6XL+TucPEwJSSkxA/6wK+flZbTTfr2xBEOgOfAK6sDbe7
N2eV1qcLJ7vN3NEHPwjwum4jRcNiJmE3We4Hl/ZdBqdwrZtAt+fNxdmyy93TexZI161Tiv/IMzCu
kia72I26Y6pe4KeeJ+FIEAXd0IFDj/suUrJNXwd8IpZfnDJM2OXGvJuhOmG3+JRwW+RHPfrWj8Yv
KUxS8/pGi9PcNp1NMit8ChLeZY6ter4FBiLGijyXgoxiCPasQtS1JTGJcjVdG4QrUmD0KfAc/jz9
n9KK7WQxs52LLioCNGdThLPcHp0D6Ru+o0pN1u4AfUXtkcXFOZlS0bLqD8hJSWCX5RPscDXE2+mL
srBq5WpohM7n6PoBBf5EuuE3BqS/dxoM4N6ZnHbq1j2/fhhF+cMhIZ8d+6SvniRYSkfYrrWTDoXe
sO3KEAXPG+CTwBCCGMdWhNFOj+ztWnIf+TijKRDoIJW9CDO+LVyIbwVOMc0nHYXUvFF7rDGyseDp
0a3i1cvXs4iApdNQxnolUY2gbsK1Vc7H3k5JPO0Ms1ZsmFB3gnI0TVz9+RBjxqG36sFzR8wph2V2
vcZxrG1j0nx6qRCndl4RfSIxzqnL+dBYZa9AitdKWjgW/gX7607bUR8m1SKOkk1B8JKIXcZ7vRe1
h5M6ap9GB+eD3xJQuOHTW5wzn+9ggC5D76KCVE7yFmZbNe6uy/sTu+kp0KQly9bJhK48f/6266ig
aWlUSNNsD2sLy+7e7yjwUclio0ZzajfTc2z7pG7+knosolQe7KxZhtiQdy5Fvj4qq9cHmfCzOgKm
dPTjRdNv8/FDsmBsHUjQNXEe0RXMYoGrRLjulxmewFudRF8nMdVQKCrlJSU4k6S8zGJVjwPiHvQY
zEK/tYcEPC/VO7Wmq4aJ4OcfSsZY2cuFeY3rsNv/+9r4Yj2I/1hvxvntlbldpZN4X/+//ktFOwwq
oLlek+A5rmZoDfsvbEWQqZK3vrXwyAjyWGc1pY3geHVjOLwTVVSEUEi5ZTaKd+D+H7wVQFJlgtWK
UHFdfthoHqWzdmQY5CABKeauMZP8vgKWv/y8SGLj7vDHTIGwUi9tuzSSfteBvzZSQvrS8VohtSdF
/8eQ5IpOBfuELusULKex1TNZDfM6OODLVpFPHMMeJAcThpxSjuTdad/1H1fPpe+eyBmMrGrPtdYQ
by9/YpWGYciTfiiOSumdae40M4yvrCWspCmW/G2Fer3OCDvseakZxjkUiampaTOT4OZ3w0nQ54ZC
NGBpLtu6x0EM+6OW4fPyDsAh2qsuYy9qmN5+oG+uxUzzeRI/COSNMFvmOmd8edUgK8ykuGkqM6cw
2qWFli/M6T5LP2a7TBazdsCfwwlfRXrppmfM0usZPYTn/VNgLk91FLY3zIRE1q02ODPN/zsaI1Jd
0fooPLqH6d/ACczcR4QW5Zsn/2E/CNxnRDt+mpTO3mUs5rdPhYN+sEjn0C6OjZCBrqkt5ymIy1lk
jqjfvof0f/48c22KV1BU4r9BJUSH17zMwolC8jO9VLKGjBDdrOldeEyE09gQwtojsFkAs4u8PLLA
n09zsf6iD2yslvOYZSYEQk3nvWgpN9SsK8LwlHjtT6yIcWqbKtrq+CqkJBtLMnRYRSMK6gJ0TAsT
oF5Pc5WeQbcjxpgX6fxm3MoRkik9Ut9r8k5ZB44l5NNv0Wq9M6dsfnT5cvtWXOyKPdymc/jVILQM
Th/KdI2gK1+WKIszMONg1Lb0mEEk3CtoqBGHyl0TMs2hSaqOfHuognZfJENlEU+pbyLmYmZS1xNy
D6wBQlT8AOTVE7yCtp4psrubbg32JPW0v3OP0D3VORZf4+yQIPjVOJg9NzCfbm43kjNBCEGzUudz
OV4qSH01wzvDKZBeNbDao3gGzAuZ2ToYiAiaB6R9EoSKyS4B1hKHJeagW7kljioe7RnnxBpPX3mJ
kodNc+k13JGNgD20UJ7mpOJ/2Cs7e7/DbxvjdxECjkV7HL88uNyJIPTeU9t4H2V/kCiU6c1ALKpH
IfhrUAqNoE70YIfrTVPTR+IA6nO1LnqO8gJWlnZoXaZAkr0/mFmRdUdFYu3VEt75QXnXM1ba/8Kg
oMn3OZDTtMOPXQzuv2tqDYqocLHJh1eomaB09WkNebBf86YeF59RizNLdTqANevIMcHElsTnm3dH
/Wv1i7oZodRnybVqiWEDlSOEvz8/a/8uYG3ltCa0W+XzfIdIsKOle1jeETEe/mdgIAYgfXiHjoKi
SE7LRTmKTcDo4qfITtdDTMBABUZDQGEWL1b+412vVoz+y7ITXMVEzLExloqYZypwnSxYU4Tr0Nrs
fnj1PNZ7izVdkadznmz8Z63kEvSAovg0EBHZVtH+XuZKgHsRWpp9kn7Uss1qJX4fWTVo0RFBBsEu
2eU/tJvjNjoJcVJwu0/N0gbiQZWL0p58fUE+WkC5WXSsx9Yl47U5/cnblSvqIWG99xK1yuGOOlKq
8o6iQ7427v8MA1LvMvEg4vwlfGjj/B0FhrmevOo3ShOQ4t31ElAt21Zkh3dR7j+ZM7Cuvk4J8ELq
KQollwyKEsJWlGMWZm60UEdBO1MrU9K/+bt7KGwWZ9brg8KV+dLDETBeyigmqbHylInLR9OxllmE
OUIzLr8FzbBFgxSfm8IUnZbRWn6fVWtGgxUxSkKHZvB6GG0eUd6Bl0zpHu5jZSSaONhkJ4s4ubvi
3/EQEtDjmg/aNF2Mp4TlMdnuGeRkF6AAUCfrSddpKcQOPiJ1Vv3MK1J7wScqTtpUx1gmoDu+m3cb
0SudWvpF0bh0FCTxw7FSu5R+paYx/rV43Zc7ow8r9UsNA4T4Hkyh29AKt9Zd02Lw9+Jl3PYdHZU8
1gx89LEylo8ZJs4smdEf5rc3kiFOIWryIK+m7slB1WksU2nw4tcBH7hwLJtbIaU17BtU7ewBe1Jo
vsjqq+de7PYAY9AVCO7NN/SPBNDxqIP1slC98CJsJXA4HlUyXALm+L45MGK/bYBbQCL1DfzfIl5S
Z7nOSTCn9728MfpKtnCLDE+z4/hmXArW7px3/cr1L34v0fhotufgMapgCEIbyv3CuAAR2u+qymlI
/jYGD6xpSAnlxSVMNaHdqVRdOIe6cXh1+NmxbuMjxBKRLdCdNbqnDuSndkNTsOK1cK6q7p5JCPmC
OLC9e9BM9pQJDn9Ofvtbw5FoGGJBeihFkq+hUHPWqQwfAoAwH2IWvJKTcRJmpcNn2ZwMfrCDpyCf
3YkOAiwL4fxf+U4XIKGlsG6lUeWxilHKnXlBsEDJRqYDqdmu3RR45W+Jd7IgVY824yM/8PYzlAEx
PzpMYD5/6fMu0qLBgjZeqrcos8QRMY0CY64fVM4cyc6Zv4VshErT2Flaa4vYkSCd76z8kL/FGaNg
oSXo6c78vrMhLH/XaRd4er6jptiDqT72DtIiIcTjwugk/pBa1bZj7VjtW27ER5vmhZFBiM0BiAMv
yfcnKo0G+B+UYKWCKyh2e+FNSSedEPbWZzWdRWCjReA3TRt2oiUCwg/8/vVg3LiHy+H28cwK2PQH
WoPaDiwfPlqyXVOIkXWgFJjj6McqeZ1McAode4/Qnlsw6Mz/6qDdx1KQ2bK55w1uujgWs84H67mo
WFnuWXVtr4ZKIc5kaqvP8nkkiPTtLTO7iStpe2TmxFyrdQx1TT5mWPZFRNxicCdPdI5y6Zo5xtf2
/si7Ezxu4n2LVKCHhkxKZUu1wnpam/0qcZdS4nKNjDAwkrnGBs4CmR3X1MdYrPZW1FX4GC1sibxM
VF/tgnV0rbnZn0U0Ghwzf7N37NO+bmQgYVmEn+ZzvyC3PH3I2lWWJV5nDdIKdYUKYYNENhdA/ZR8
243hZm0BiZLY7rzwQybhv1lrUE7AssTc+c27aWEUQHW/urN/em8jROVMwfSy7tzNMnOPLbwBqyT9
mXDm9Rwd7MDwxd3df+vICcY7gmxPcZD690J4CA5nHgEMjzdi2N8UIulRb8DiNrtJ2g/PhNv2OP4V
DD2eTy90i9vfZtFvl0g9ZxW01kZqZ0g9i+iI4oMYmXtRoVnZbuHQi/kuxaS6W/FF10n0hKI61Jrb
faQ7aRLtkWeD+6VAYqPPyOjY8Wxl91CmSZcDdiQm8KmZFfsOhLHZucP+l/hazAUJrj1u/eoCAc+M
x31jtQyUMmzJQWP2Hjz8oxL3J+GbNHliHXDwetFdE4XyyzfzSpK7xX/fG2dM1x351XXjkQ0HJq8q
ueXYZZKeeDcY32ELehm9WFzeh1/alHImRNPJiUo2e56sOEpNArXFv7Lonv8BRN+/48ce7r6mthAb
OLpB7LcWozcSQj2pzncHbIkz6tWWRjLBoFU9sfMsk5r9LSbAPJpF30oDuQMrKP9bHqeorvu95dcG
qtbcBe+hOCDzHaGxEN5C6clrChBXHcaAN52j5qZ9JmHFD10BpfBs1gRj5yZzGbMzsSbI9KHKW77l
wuwQlkWm+no0y/G79kmDFQv/b/wjTGbzQn99YuqYdg5lnNKb+Iv3XbFR5/o611UbZiaGBzPc2IzJ
dU+s0tTfolmdmL+vM7qbTiCwSU45pfeBGMJH6aEuNCPwgqb/vmfTSA3pDq2XfACcsQIPLWnRGE3/
juxfm9P1ui/t+X4QQ20mNkwFU9ddg9lhuyQTkGgM3IWf8C9QIROH5YraHREQH29CH0yZ/Nnwyrjv
JkuksGV4rPWyf5XzlabQ0D09yFdkTIaoqFBXwVNXCP8Ktu/QMHxOLn6nYMYGgoKra6y8Ce4YKOkb
Cw9o5fNYz+BL8jr4JxUSqRmQ594Hm7E6BtB57GKUGIjZG1NyWFoeA0N3yPTMO67UTA/Xt18/Kmjg
s9UrU2dEvbVs2HYualk21LEW4PJFQ3fgz5Y2DbeNW2duVK41BTLYMiNVVf+bQ6iYJh9I4m8G5B53
8BZ/uk+CO2d/Z7LYurlIqeZtpcqzQ8kRSnwjPPnt9KfNmd6XpKavzXriJF9eJn0JCMjkVNvx/5FA
isMvVwMmdngDQppiSABoWJ3+4s7kE7QhZ8S+984hRKlV51tzhOLhckCOGO2mSIRYmb0fgRz/nsLL
N+16jc35fY5LwvLFs8iPwV9DfEBW7mboGyr7NazNUCmd52TyomoIT2MePVzoU7fuGKSPGh0qbIym
ehmLiSYh5dlEL7JSPG7VWbEyDuM2gU85C9/XRAgTNskxfMMU1OFI/Wb9iiL3wDtg4YxyuXcogA3m
VwRp4ka9zUT3Za9Xbh5bhc/G1hgq4cloxGKvL/8MSloGLcdAjmO9Z3tDHsnkMTJ7fd5EPGrtvcvb
+QvaJjAvofg/flSBbcdIPCpjqctwWDf1iGm0DIw6Mdtne1v81yhkDGMoSiBWHLZE+0MLBXTYm0xp
+iGfjsZBHK/diMUf0CsZCBZ1/ZPEed4GPjDtBOA/4CL1ugDNgdjufjEu1jsUA4OP8zpRpPpYh2DC
y9kL0Q2GjO/FDleO/LQNw6l6o6LtkQDArzeik7iTYzOw2B29nUWs2VZ+dbYmwPO/zligStUlz28V
n/NYrI9fpw3R20gPbhy+f8MV8GjDF+sG40Lho6jg7Kwh6xXV4pV1OEJDzdf6OBtaei1mRDdNuE22
yeWiDDKedPg860ZPiPvCS5sZiL3a1+RzYMi09uiIGueJjfjdxWyfk9yAEE1Cp1y+i4y3h0tTaiUO
TOhZY1Sst7PCbGntBE4FOzpHa92th1JlND0ECgwK39RJce4Ce6bp7XyvUXvy2Ku7qaU0SGD1ht2S
Q2JshnyAc2W5Or2mA7bolUOKdFhv+tco5oT9KCzRwzrarRo3qszBv/LO0h34nf1nTThqD34NkuuD
za/3vJ/aX6oGJu8dPR7gjeRyhmvRktDVz9iujc7CH4hnyk7wn5lIOYCKPFX1VC6yZPpFCtrIDYw5
8pXNpMKse2y9B4ant2wJ8ATnp6pkKweDUAN+znGH4kfG/QDrNQxUZNIi1kFv923CaetTs0lvLmzv
KEeXo0MWODSesuJcZUYqheC3Sj1zqEmAfll5f7/uWMgW5xG3JIEMcG1FXazMa5tjinnKp4l1dkD7
4Ko2e0y6vLkq+DU8ivNqT0srvrpi2Yle4Jr6oobgWpAszFS9+NgXS78ve9/nfgxvl9Yfu7fDpYOE
Zr6EolVOUc381p1mBlZgtLRktc+VCYUEy9KsbSZxszyxIym2ZW2zuTSId0ubCtRrDkN87kT7Im6i
xO8qP33W6veZbuXL/+6c0PNpkgzTLF9T0fONzGnVmEIJolvLQ0ZDxkK9TaslUSAF0m4EFUAMKXdL
eIsb1C48+8H+rp5kYEgsD/lk5gy4/65psrAn41E+1odqFsqySvC94+AFHCgALxRRmLU9yd9vlCv4
qWxlwi4zQKOMl5hfVyPcbE+RHULbmnG1NiG88ZKgux/2/GZgmLsVdqjHcPrS4uG3Qrv1hKpT5Rzh
2itzaDMg0kVr5QCkUhT7rqN3FAsjS3UZLY/i0h125tsPsl3fbapT0BC6u+pY3kaYniCY5y2BiL8h
pkHx6qfISk/PTUa5V5Fnf8fq5UVc/cwAsrhEOa1arydW3pmGg9YYdZJ36ni63CMVpqZ45SkZ6xer
qMjscJ0i3PnzDWTC544t5gywbOCvObdryyX3mceNUU/vNDu3WSqhA7scqW/9j8sYEwkIo4naRMau
lohecV92h2moDVwfgXuqpD2Vm3HeezjkJyKbLGSmz4cloS5KtlPuQxUKdgjGGuC5jjnTfKY/Fdaz
5iflbKdNGWjQfAWfK9fZ9qxhrfuCblY8jDO/u8FjI+7umZXqqDjAjsMiTdPRNxE9oetqksNYKeFH
VaEl/+Mh/XmOI+AGm6d9tuoRSe504rm9Wr0EcvrgbfMOev/6lgsx/+TlN9t5IiNC+xqfsgBlPf86
n0jNC0HqDolB0UyWm5Ri4KtNk+02C61Ya2Bo+RSesPVh0Yp2EmFnbqaYd1Ztykt8/VF4/lXdXhwf
3OoLAWCDnkY9nQV11ytiZQSVgLcetfrA9a3szgSWYufWxb7oTIdA3wWbXca91uQxPZBi39BzEUhI
ZwQt2ST9kGZcploSYPTXeQdYEr2fSLosMoh/ur0ASShFEBbbo5ZrOrv9uTzNS4pxFxvNdCRHa9TF
yvvNf42GNFBODTaectdxQ/z2r+2xmkFsX6BDc6kkaDS+sbDnvPi09PLDLnLAa+yh0pjmQlFNTFES
ajdta0xlDWHNDplnnoEgGoJTvoD5JrX0XkygtohQRA1lWq+N3JXA5V0mGAp7QrURatiNriE0Er4k
hWpE1Am/w1nI3cd8YG2eP7xnaPwXSYwUvlpxHYJvHMo7ZVhht8WSxEcxSL/KVzHcgO8UoHw0m3jM
YYUMY6J/CcFxNRimNOpA7eCI+yl8Vtuhy53DMThOXhJYGhHVnMgOs+zaJPfzcoyPs2ONWbyyfCiq
tfWZpz3KZlwhJ7OeokQbsQRV0Xl4D2eJocm/zz2607jijS+MX7Um4052QAl2N1/TBqVtI6gcf/82
r46YwANzF4uk7VMg4qztdfNBl469p6TrmoEMA8/f4SqqXNe6J2AAYFWPkB25KMZ4pS3GohMG2dCB
6mZB98Xq/eHyhR5XPPlbmuxDQUtyOI69MG1YCfwA6bx1QAwZl6fXeYNfEdtBSRvXSxE6AGyi2Mwg
htr9m3FpeDBLEqbsslk5cPNMKNVKByNZa8vZwE6YgdaTpvER5hikiDrRZAJqH9GCzQmD/G0O2yC7
5m1O5SNCUAe8td5+w3ufVYLkG65fY0tqueEKESCOwksNBLm5ty2KykoLPkGAJ2Dh4w/QNMhCaJ6a
tTan5a1tT8vnaYjZS9mKRURth8YwzjXkdKpURzlh7jWvuVrC7kRGKYMZcmNXbwOd5nfo8zo3HtuW
OMWr5SnFr0DXgOi8wA5E+T6f9T/iB9V4v39/zsnE9tGHTrFWB7JBW9MFjlFmBdTO6F6uUzJISSG0
xHl7Kp56LSz5uo0g1vT0be9CCi6gEfQSoq+FpNTrLXDSjfBMjVXAXZnyrV63Pn1l+KZwSo/LDcy0
cVzzDWOcfiNybxPSfWbQ/5KabiuVmXLsX8MO7UFCqrg1QYrqxGE9Fk3HfXpP10jVcwaHcKeSvZC6
ibgF7pVJg8P+KTh6eFUMavX+oj+FI3pLtqnbkNEsfG0qP30KrwUaE9xKJ6/XSRVzhS579ILl3eNO
sXVvbhuyYxAR4gOjrvv10dN84SG4BhZW8/yVvySI52oe3kYQ3HRNXy6TohBa3f462ioZfDmLD1h9
yuL9TBNDtNVQlh/VJ0UZmPWcHV9FobB9Loqz97T4IxDKEYl8mNQHxtZWuTw5PKIOY7xwMaPabGBW
ncSFgE/VtkiliAf2n+f2/ast5sSZrfi9CnFacyotSxsbIBTps8htVyOK2UQGcNc3shAdLJiny8cP
XQUtDWR4EiMfeVEOI3OcV8G4ugtM6z6qeTi4PJn7vNUB8W8TeK4i8FG9zNgkL6+HavkcvS/l34qB
UH8pfGNBbbLmiOxWIGM/m3k7bBGm4xrm5HR298cYtGnmr2HpJQiwNNEYt7/Y8MziQYpsBJ71CKD5
dkfuZvF75R3IDXEbtsNcdhyQxsc+YZZmJecc/fMtSlaEQLliaYPZJ0XKTG7ArCdSXaUKsGr5NTwE
08QEnDNlah+SmwiSj6fGLKK2BDszO4urWX/WtsZJbcNPfzVhiHELdKwABiaxq6oDBr/Q4IagofFw
6Qc2XhROILrytMrC9NllW9tZj1wsk77Fu2CNp6ipoS/F3nPEPjZfFzd70Dr6JbTmYd3sZrtKyLNI
bokMmEXJqe/IPikDrpyKs0TzmG5JRKhZ9ATgjGD1gFs5zOgL7NYVJ6DhzIMcXrwLhXW6YR1gJ8T6
f/vQrc2bmbeamzl0eboPypCdGNYhVqBAJgRTmgQtx1dl9L8Lj4c9N2YJVaDJSy5JoZ7lD7hAKf3x
wpf9QF8vgUZS9dpziGeG4rUEjb7dGhdyJAyVcJXfN/Feq4Ksv+RoAvpMJRlLNQq3zWvt0qgltrHR
iARGZcfxLlU796qWIjRXjPARSNjtceOwHxSlkW32ItOpAMDRkDIsWvteG1O6JcP2jt1aFC3cWFs7
dH+QORsHVlun+V+ZMJkH839JTOQJE8DEpw1sJzv40cseaMCRqL2ddZf0tU2xfl5M1B3uSsg3rUA0
vNwvna703Au+9imrz08Ee7LvpoIbSZfRathTpufUiFSBu/MRAoBtrArcKXpaEx5JxhcSHJt2LjWK
LS5+xmw6xf3XOlZO+r/R16aDluxJcTnJN8D6xIUE2U7XO8LvN8k1zvHpW9ZeM3T6IlFXLlzHyo6G
W+bYGjoSQ9/dbEyza+y3En1/PrjiHvHSYHB1/uGdTzAt3PflXu8S8w8kRWRNuaSemVAGE4LVoJ+R
MR75JDRfdprNpGInp7fyQ/1RmpJFwn2ASX/kGpXZZk63JUGb6/SCCHrjJ+NyP21ZJ1QyMWqUF2Px
wQp6ULYcgPt1GBB/vb2wuiEFJpFXaqWDV+M+IQWU2gQvbo9hW428nAsqTWIMqQMZnaXlHaxMemdz
2FEamqLZJON3roBkcRgc7rYcyv9cNx0e8WBAdZtdIE9VGB39gcj8BJxNXyuNMYo3O4lEGx+x6ThY
HT34BW99EE92aq6/Hj0vTw4n7cShmKWEi1x7JCnPox+jDRgBcOmw0YhxoInUB0qf6PXhfjlG38E+
sP3aEZcU0jBaOMlmGkCWuL76ByZVCr8TXvZj0rVO1J1ceOdJcIqfV9beEbKnP8u0l4QA7vCN5aBd
nHpUlN8z9U1+D7suSOqG6v8XK+AZqiJbbjm2lSVVj5PQJRscQMC9JiWJLXW7eAlFxwDJaoCs7Xbv
EvibhLzTCbisUrOVAKIYOA+3fy1thugzFT7R4DZxAplYDyH9kUTDuYgEj9K6TZgsRjnmJg/swuSO
EYDbJ9TRtd876homuxsWjHC041RNQbKc85JQj/Gu+wkKuF4bNGfXcN/WPZknW9u2Q3I8+hGzJOJh
9eOzsr0i/qfPtRiC56OXb/mLYXCmu92TMhdU2CYeBNHn81inqF0uGhE2+DDSTO4pnPSmzt+LMkTH
qzckYXqswtTsMZ2Fvfl0Wl9V5eDBwh9XTRI7lFtOwYkYzJewlBXUDAlNn8UWEyPqX+Q6J92uPsmA
x6bgbqr8kin71EKePA62jMHGMy8356A/tXT01OeNL6rR/4UCzzVQM3D6XmpdOHeXuzPdXD86ium3
5YzDXtyqDfMsigOFxujV7RTVdKFB1UtEhOfokEKIm4uPV/qwTwJURoYDzQecXOyW8tTIR03DuppB
N48ba/GH2SLqKupyyeOSjL1arSsJVRF5AuAVPNsPYj5yI+XjkJurXT0aVJVcUy4L9pQ0wy1/u0md
vmmR2eYMkNcqJPrYVW0e9A5TB5BJC3llEIwWpKgaFaMIBHAPEaWGv3fHYk7uNe56V1AhXpYIIIXg
BL7OVqAbUUHGE6WnsbBmp8ZOjK5X+eLZnogaEu7rr8rQP/y38qUOaY46AvakccK5vpCbHc91/EUO
o1U8rGGSG1l176y2Jh/sj5YimLtJHViPNL6iBELns8ciIKwR5UMnPydZk69ek/P3rvNVKTGfG7Fm
E358ZyyduZSYRS4gxI6GVRwiUnmJrFy/k76S84mh3t6QM6uZW3+1QYWUEhbUSEOcoRDoDTNgklf4
5gXJ1i9iY3WRYxfBqgQWC5oeP+whXQUTdLwfh9QxNSvGHSjnWE7aXnuxdwUqsCb1L8x6a2p6NnQL
pz8E31xOQkdHvJ6kO8/7SJp5SrFETGusVd7bfwb2dt3WEpshYqyh6jUUD6071r+lcxByS1f58PlJ
8qfLIre1jYo9zgGs+3bGOGA5xgJFJXUGwhPnf7Z1R6d6yYu1CVIdL2jQgTbub51MmNAyrhfrbH+T
htWIFGmsojCVInNfIPpqAosBnveQ1NEPphH+k4kP1jaS9CD+YEgroctQMMtxfXqNmtKUsG+ZbtcH
FKu5MypoKu5Lklo38zJg5UAs/bpnKhXnFBOOGrbNgUnmpWfx0i3W2/jreyRk+x8nN16h2nlLAlnr
9C8xGT8fQhj+Hrz5pOkj7f7b1p2PeVr77khFGDAX2j248Tl4R/m/oQDSSiErWMHlgJ426xPSz45X
nQLcOiFPGdnYwRMp6odKS7HtKJI+/ekKHcLzpJaH1cPAJ64EE3DTjROQw4KGJHP7ACIkkqV3QvT8
8HPU4pao9E+sDu5zSsWDmFyDZkdz3dYHwHJpTaS2ENz5twhS/0JQWzF/Mm1J9mZqtIl2s0BXebay
lthpRsUJUY3Loi3fTDWoddtkK2Q+geC0ff8QX25BpjgQ43dmqyEQH/RaAwSmDSZpnGO/AMsRagXw
O2Sy6QxWz+QAGlK/amGHqcabgFyQzZofyLxafQpXAggcWmVN3aF8DHsbE4HoR0n7uiESqjim0XGj
E7Xfn1PMOuKkYmCAvR6puKxA96Asj+mB7NXmhaRM8cBWJ66Ja8sndOSKlfH35vv7IhyLjdGyUAx1
iq00w8+pc6De3pKfQS9/6WvUye1ZEUQ/zUO0yg3IBQW3DrbdJpoi5Gh/SUyWC2qTXBPeAZY5Dv5s
EaFqsRF1z374yDhG9VMSAT8yImJPRf1HD1D2PcOht23URQDrfQBl4zdZjfkPFFWygtNxpFmn7dmR
/tm8jnU8w5xVmEMtMXVbhFUfoCcUAa3AfmRvxr598s4BDYpVBDd5En3SKN0f7Bgl6eyxYwUSk/Tx
ao0hYwfEF2Bz4X0kpIVt9tBWrEJnzJLNxun7lr59nmwDunkgBL2NmDpgdJQqjzo7HWjWTqxZGKUn
Or2607YefJ6YbjuS7W5r7uKYfqY/wjpQw04wyvaQ+vNHj2m7+Lp5mpzb7w3yCGZJY3tTpNObmYQN
3pSHVbqmHWkWAcNTCsdXIHdHZcmcCdZ4WPKxcnC+wYp1yh9B/LaZwIEQpc5XHhsr7TkFFzlH+iwk
+m0eREco4/BnL5grkVW8ZywoxlwNNYekGrz3FttsGnh/pNzXazXQh1yehmgYOBeZyyyLVB/+Ytsg
WnboshwcI8E1CRyXcR7yHBwWWvo/z1Tl1CDf6JhD4H9u8MI1wyApS5TCEF3JuqBHJl9yc2wJZWj/
ug1D1S9pm3D6JowxnrT8w6Z50K2Pq3M+D1ktG8zipbOkcn/SOusMgL75ud0uz/afnXURyL9eF009
zjl0KWCLCBind/05lQCMy7130F1aQu9doQyJ1AoTZZowNuEmxxaBTYub0LH6VA7bQZ8uRMbcjpi9
YQcW54mG4AT4K4XXZHcLfgTvZ+yE26MmqH+DomIZcqdGiqwuKq6XXkqNbN6EnquX0S6K0yVT9Z4+
7HX2eeINh+4evE8Cukv6bfuVzpGozA57aByNBeIRCJmXvYdLm2nNzE0zgrQA/hWGuij3wCc2krEf
bVbvV5aLET4vimQ3BAozt+o2rBbD0Q5GL00k3HzdwOcxv+uO5ielTkVmrOA9L++0nPvpLNtWnAFX
O2JRhugdwUj0FhE7GRgRearqDQ4O58I5ye2sB2fveKUZaOlqJT4yIU8k6FzbygNzwoXRQPxIfFa3
tuGRfz6zAPQZ6dmfi9sCLPO4f+A/rw65mouNIQnIsalUH9VJESAFKRCvvwInK++6tFG1/+Wa6ZJI
6LAQEIeK67VmDFt/sA/NOoelvYtzZjffVHaHN2ef9VzsiAYUh29GWbbeTpViU/d9PbC4L+1BqU2T
luRljYkvf+AFmxL+ADk1NQfCVzp/GaYOnMJrXMKqJ7CxYwvHEoHFqmFvxUq0LxOosqAj9GXZJhZS
8H8dI2Lp6vaWPaCvfFoEpve+dvM8SVnBDZKeK7v1dXLYhnMWiB5hmDh5yH1pr1/rwZYYnliCfHjr
sWDHsIi+2uAitEdGok8o2ip0/JGMbID2OlCnzNUltbgDscx6uj9rj0KP9FgqzHF3JW5ZigIaJDgR
dwL5qgFOXWKUhSkNp8sV9a3eTbdNDPfN/xljtPpvjWDHvlDLIanNng6VTvt3iVYErep1k2+iSdVj
i4Jhq2PfaxwfMDgr11HwYqJr+W1QGJHyyEZ5g8PDychyRCfBx6xn586be+yquEw/ZKjJAww8Uujk
f3W3UsncDzAYuCzxEqibBngNt1Zbvd41Y67eNaK5KW/GRnOTW78F4zKS5zTZyjj9Gr33umxDTExA
ShK68JbEG//aDIqu/Q+MoToqYvejmBf4rMNmmHQpzbrjUDQIWtcSvli9PDwapHsyXTadkI6F94iP
yK3HtBbF46sukXGS9+ZLUBMc8Jidwn2elZdRDl3k6OZCmVufZPG45YkfYl+ni8JQpqmuk910n9rD
JvD0cHzHLrXI9Z5zLvruacL7lw6Dnc6Amv+F8pXCj/v6eg/dz8ymV8wei97l3m2S3G5hrLitb0z2
/sVTlOn9lpHELmPBva1SvRGNm1WJ71Drh6UW+N0ZhdJ5Ymty+KAQqD/OD72m6J7GH7vZnMtCyTkL
WdlEuniTPVM5vPOOW4d6O1+3tdggxM9cMfq5omcXU072RxEbAyXSu1ZNH44tFme6qcJ6OXOYBYgW
7LWpr1q7UKtAGWqvqLu5m6qyBFD2671GRUUncHUTK4pNMxbEC8oumAoBaB5tfSdTCFB+UKUVVzUa
Lost+kU/rvhW1UR6CIOxvm02ayOssBf4JiyrH0v7J9gnxbgD/jA1EHlZdSkHPfDD3x91YvdpALFt
euLO2SOcIMp60PYhe2C2uHIH/3Db9Yh98ah+GlhMx+I4xSYuNeWJt1rdODTiV5q1jSHrkiu6f2n/
E7uJLYnoNGAr0Y9icjjiQWZJZz+6OUXHCHlOCTee58G8lQ2HgLVrdFF+vTEPG8C+0c0RRUVE2gJK
uoaAhmUHaPvdkAZ4ds6KsU5TvRnR0fjQ3k79K0yoo1getIz1n3FFh7U7B7r1nEaZPsZ3NRnRKXKV
TyyicxWolbl6dk7fu0OIYH/UnNozO5vnsQBk+ET7U59Y3kX7XBGViGu+fIZCdOfFd20K1bN4jv4o
FXyOeoSYfDgdXMaacq1dBlLEUSA2dfHiYN86vcVBr7VdPlUVbdeEtDXEl7n2kNjPW2xjSDAxTwBV
CJkBSKAx05WzQqEZFSLhEnFRpWgUuBkucpAH38dSNYMoK7H25pVYlbzmUejU4X9rlRlSSGNYooN4
UdUUSvFluj6sOTa3vIcc4GmtCPHsH9juvhMwocuidf/r2906bYN1Wr/F6+pjsuS9N2COfqK4QSaW
CP1EHfwzoHY5uiuALM6kqEzj+Pae/3VwCeufaZALtkr+6m9Zt0HZvZ2mNeNStpSw1xCA4mVnoo76
GZK7Uyc5XMFQaK0MSDlacKTadgDjsiZ7MQRCGaelwuAZCu6OgICw3Fq4fAmPz6sVwIQ95THlGBat
qMGt7G9pJwtaNKji6o96MejjK+GwAdt3rMtn4uNwJk/8qTeVCgHy1ckbFor9b43afqfsM2RN4Va8
zSD0HEWu7OSGzVRk0/owLHuEX05+u1+R0sIwRx4N3RVXyvdKvw7K8V9DF4Eeqh5ka9Kkrqcr+4uL
6hW8GFnU/gLxUSgvGBjig3PgaOK2xxepBdYOaN+2GcNcllUyP6tJey8ThNO0xh78yk5Za0VFy0p4
qipmyQgFJMIKuiWr0menRFuNx41t6hMUH3Ed3X+2Q59EDgf8ziZSrnwrHKcsukNOg5sT1FBwnTwX
nrEQusMfGWPsCmt2QYQezbPgl/yeyQEiLSOIbDVQNLu8M6nVpWh6W5wK9CEgnZ4YdNyPPwLoL1q0
cyQXw6Kf6otr/O7Xhc/ijLaeAcEhoabZTmjgZnU317X8U+V1Rmo+apy+5rHSfwcC2dD6hUrqAi+v
2YD8tTcOVkUHVjvZgSXdEJ08kCtRmjXJNi82tkHDUMpaqIJywBvWyZOSkQWetudLuilos81bnm0/
vAc9Q0qYVelntPmowcmn1S32tTcvrAnmMNURTs7ekF7iqrhhNXGvgubV3hFzEIsr/w4x+ht2qGNe
Mp1g+OLtFjbyYEZ2x5hT6myjSZer4A65Tw7Lu29cv6OovkZU8/GtYPs1b7USVtFLgXBZvWuuFgds
o3j+V0CfnCzQZwyfE9pZpjCxhjoUvISUAnryRhb9FFIJLhevAUaSvFVnfF47aP8H0gpFdXQ86+oz
GKBSyAYsaIc0qBiS/0GEi4aS1QIaaTspVx+qlsH+kRF2Yq10SwSLlygBdwTSd6NV3Hmxr1ZfpJkK
UeIVOD25TsE9l1iLdjev9EtPrNnITWdfl+g/HtB5MmovToC6kG90lwcq67RnUAt3xSP0O/D6dkWN
FF2GVoJDPWjntK2krr2kw1C+TnzKSmYIn7gNZnMzuqi3tLH+pYPKLnP4RTlZ4VEB+uVcSU2Fe14V
0ZzczdPE8CCC59SRK//4tAYUYanYjnEmM86Guvrrq1ouK1SqOD3M5YUQ2vjGghqvCjXEb67F2CpU
xNItI+v0EkUOG7Sb/YIUCcsmv1McaGH9z8PWhebbWallRY3v9jIW329JJxYTutyvy8JwB7J4zA8W
zENXBTNarykBwiPpHU68v49B3W9hkbmwEvHRNeWSMJm/LHuYq94NzbrFW3x0MTWsQvldNvRLVFDG
h8fE6eG9MgyU/rKAwKRNnEX4JaDpg5k57++YU/frFUFQu48OhWHzQ/bbSL2qdcJSvyU4foCuMTb1
QGRXF1H592ggpeeMmqdEhTffFZqH+b6c8W5Lc1uHnqfSFILDxewMnee/Jymzk5OxcSwuDvqM0uVS
OwF0WzaIkmwBFsWj8Y+B/UmVr7/1i6BIOTDrAmaIvKUOXXg+LpQFB1TFGCHqxlBsr0Hjk2ztVJeW
ZUxXUZ1/Du/Wj1E5EMYxtbrb9kOLWUJiLlFwiVeyzynjRV4pmnhuZRIVQN6m3I1ELWSoYF/Ctzx2
B+yh3L9+WfHlPpWw1NBg0F00Xh/3J/3go3Wp+yaUTp75wyivGswkzdBkZi0by7r9fKs0ak1WeLUK
hy6rZLJQhNSEME50xbA7djAqu418RdfYMKRPUixkNSI4BwEHX34l8+OFeZCFXvUqqAbrfDOrQPlt
ivoyEX+LvrhKOwq56r4z9kZSXVub0Il0pUoUigxdCOUc9zKUNtyl1Vdm1H5v+pHcm9uMgfmbgCGi
5TC7cbn/KHZ/TthGzhrjCFrPTkSzwWhp418ZbCJvOIt0dSU0R4B+x2sQQQUEMePG3R/3wRjaHksI
3mH2nDWGO8/7Hbo2/yCmIabloqog8L6ZPcLqqGeAuXrRVhcZ7LOSV2j16+UPuWGXBtmBN/iPerr9
tOB3NqaCMrKfcjuyt7f3GYRup/4GYh/1Ke9ogrPXTASNuFp8gdR4YNfH4dE9TohedHfeghoBa2Vx
t39CyQQCgTA9lXdIp5msEA0oZVgp4qPFgRRLu6YTfNamMaMraMRlQh2KjaPm0iT4/X4PMCu06E8M
eXR3t2Rplqavt6L4eLv7Lm0oNGkccEUEjwYsRoztsNKLLdr6JxrYL474k85UNOdqU+LCt3hnWSaa
JOljBnUG5DBdK+dHxfvNMz6uLLMWP4PQBSfZJ4EBhlaYnfNDrGW+Akk7+wgVvNv0tuBNARhOHsu/
6owzyypZ+1zg+TDtqbTren4zHRYvF/udbphG9KVkd2kl1DAH/sE7bxWDr5d0wkzYvcOTSAlG6XJb
0ymhBHZn6kzqLJLwZnM9Pl7Rw/bEn4qnI82UpWcVRhx9MPt+PsE2BxewacLdZbDf1n1caEjT8WYg
YEj4Xi1D4loPnwAOxdmPnxCniqUGWT48DqLg94JA4CqHUxsK2jsanJkLhYv7A/7Z381O37Bxy5j0
5kHCrA8iGiIh0ck9jFp4y7AdcFHody+pR1SPfRC2P+IYINtetJzqQObULrlnNS8QSJoZMd355lBf
8PUxe4mhCNUyB8IUBFghLG4BI/rHY11EljhHasNCTrfRi8eo7M4VkP53l8U+f4ZrF9u+CtzWns9a
mEIEqL0qC8Gi9j/MuVqxREP3Nq1Bff9uD1y6sbV0OqyBjFbsf4vnxw5wTAaSPAr6LENwO6vPiSzu
79YOijaBXYRYkmmFbEAjjJUtLD+L3XUAmgQ0hTqoVwsOoYgnWC9ESY9VLsy07I7wzk5J3PdOEXGB
LMWRcnOOOz5EB2ICtVZjrBSZUISfmtYgcqEX1ZabkxABXnegOZ1iEmAJvJVb9ivLtdwr4ebskFIJ
GxWxkaBNZaqBJmw26E4R5I9ubSvOB0F84Ev9R1OUxrUVeq58mI54ev5eTgEA+N3cX4KJkexKaQlN
nLJgejARLFa/ig+JUb5Dr/HLfV+oAxHenCIhQ9TONfVhD0nRsQyANb1ShLMQIfOeZppkV5xbU1sD
g0ybaurdRRBFhzbneBNvSI4LbwNuFM3L5CZoxVxCcUmsF5dZSQ6AC05I/zDiGAxzWrOJ19xtSUjM
DVn5vQqTxMcI/qKmAqlr44nmEYDQlcdicI+2aINaDCctDdTdpi+v09Vdwr+WoCaxUtMtlQA4ncfE
OkQVX5NK+gXDSqRWAkNxph6mVeZhgqcBi+qpMbsd0VXN+Hb8vGa8fs6BVtk5o1+NBcy/YA96ipsp
2+nA9SJuV9j1CYkJNYNr7EUnFsADxw1FQq0KYD+6WKakCA9zg4vRSOsAM9hrriKhC9I80n0uFTn8
yYuUYu4T0Uq8XrelLbmAI8mV8FQWiE3N/zGP3tCRP3gFtdFR3/OzcXDmbl2PAHC3c7mdJibFN+ix
0hj9gLeVHvCzFBZJ+Uge+u0PhFkgOLPelLI1giMGWVfZEL7GkRW0Lniti/4l7uenCVJqc+frKB7N
ER03OO8b8nvpWVw808nUUFnJPAthEgCcaGfMOL7vFNwCN1HvGsaaGm7scabquI86KB/XDiM1jfM8
C+S/RNDmsHAz2X7ClAWO5e8+NcO3mRzA3VATITe1hTRpy4MU17yk3Ulv+MKZdEFX2sO3mDBZqmXp
OGQkKBVO28ZJx6WhEsonVKZL2ODrKexooauoFFDe95bqSJv03gg1ht17AfOgOE5tFleD6v2fFUXO
4XQkLtrg5GlCGByXm7VgMt1rMs/WeEqX1fVz/y542NW4LV1epmuYbMFGFsIp1aelyQqzRL83Gnm3
P/S65HgRbaTrWCzsHOlq1STBHYPK2Qdhbksj4E8Ow6OTTqU2M/WYioAP+mV1i8Ayf0FsXWoeay/O
wTxNBCvY/JmZT45s8FTKo0juTfv0mP+M6XWcmQPnD+A5t8A/Q8tz7no+SCOUZtQhZaEvboOWdBWG
uQSsrD3yOhP4BkZN3YeVSjL/msdo9We5xiQIHgkG0eJCrO6qPmTb2DbA/36GlANQoGajbfqxrmBM
TtaxGv1FqUVo4BBUfN84HRQan9RW4N2vqGPW6zwj4cJIzevn0BUc86DUpBDk8ZVhFImLYXZk3RtU
pwCIcLswRSBzI1THCA6iAo7IebJl2YBt8tSgGDOjHFwOpvtspB9eZ9v+A39gLer7UFaMPelMTYHE
z3V/3Gaz8+DZRYPPbTwKVZhVrStsbIIRtAhiNX0hSun6wcAHlN3zEZJPsYlzklRVRN6qNQU/fF95
98pxAK9Fc9Z6FlnsNFUnxbeYOiSsXyZKCHgPmFNDUjoenDQSE2frQaAuFqpjinf2IvTIt5aaIw88
FWaioeRP9pJgY8Ldr7VsutTo8dRJGixk+oKz3TdFtT1N0oZjOE3dpVTNM058WdDEMLNEIYNhQuNF
MJsvpaX8mnrhwO2a68dVkR+hlEsI9+SsCDbuRGN3f+uk07VQYaw8+2lRAKZqo5ffAKZKsu27wizI
R5IRNKtbGccZvoC/DJZlNTdP1VuAnfcuXfUnvGG4tLz6hdEYxRWguMSiifimcTXL+d7JJzyYoFGq
1udQ+gbyjOTtuwH/yaW0l/oZEcfpDgV8W2ucyds6lXZ/W41EJ5phCHp0mPImah+wm0YGMgFObaFR
XDvYBMvqD0JnHkdmN0JkbKN9m7gM6rqsAmBOpQb4DO6BF7+X04EOoIROVIkU3QfK6aWvcPvgoLzK
Avdj/gKsZpfJQcd4OYCxPNod5XxA5ueey4G1bC7OlOkMXdG9ImLDHS4FSwPWh6CSMXKd1dgwBRGX
nnKJIDJ5E+MHGYfTBF6fD5YIIuOs6kzHqzfmnO0cHPIyEIRQtiatnis+RAeUcEk9dutPcFzHpls8
BISqOz0JJXikiKROufxpqFqMWfah0vrtY+IX0K1bsGNmKhFNP40UDCqoDq97BCjUsd2Z0hy/lsAv
WEiHAappX85Bm4iG+LEbiJzKj5DymB3lUaQs3WIOxJSk90y1WF/Vtd4kLfSYco/OCS3v86JrUCUz
vTkDRdfxsVuR7uq7OSzoC9wFiuY9AgtyA/kPP9QbHAg9qYpDjKYEZG78tD/hS4XKhRlT957VeB03
DeOiMF5uVhheS2g/NU6uX52TBuSV8KzwbOjJeT38tnrERuaOYifPNxivx6bcsPc2+pFee/CEWdq3
ESVYDWtQnLu/G1uemGLtl9zMIZCvsOc8Lmqdfg9s4uK6eDFM5ONeTLwGR56eNASU+Qr2lSqO3uka
uuWVVvC6jzHKI+HmlM8kq98Ej6JLjdOyEpBQWek2fiK4LhcC3Fbz41HTVzFsETGmtvyTxV1Ylysc
WLkMWRltL87oOLZMH9JZTGcsbIidSvjqbE3ATIgEtcIcwYuhuphDUTl8Tc4iDNaiOjVGb6//BJaN
US7xEmNkHA5TvxEWnVNbCQw6VbVKHUeGTcM+tDzuNITReJ0FEUfZbRGcaTLyofF9K2SC/Ig7LcrG
b47sh5d0B/c++jhu4kcVUSDcylSVAUga3gxn1OC8+reAH5Ck4HPLuIpV+9I8dqMwG13mvNjUYokV
eG+tODH7wAkNeQ1VtnjzmtSbipEG6pAOEZAwGqZf/1zFUNKnRWSHO+lkYZQ+wdFiXjwtLEpbqXye
/9IzJxztw19RExS74SIqSUN0JH1uYVW6n7LCTA+1X1txVMnmbfe9mbQT5UBEiP9irSsDwAPAPAUU
SaYsvkYAAI5LXPwQra9qy28C4yATuAXkM4IsNtH4/Z+X3CnCz0DbOB2YrjbjJtUvC/+Yh/hSjT2r
/UpUaAF28bAbKOhcqoD1OzVOSTGfiZE4Ikk5MnvCS1snthcd6vM1+HMtNk9Nigvinf6bspyrRreH
zLoZyrNowiLcN9lVqxZquKLtLj3n48aTpAWxHmcfAKP1iIyzX/cs29u4UF0vV2B+bj/Cf4j90ez7
5PW8Rr27F7FzU1zshBzltzCEQGtHn4arp1l8Tfi3tVHcyeVejnXOBBGWll2RRVohZtu9q8M5cGPj
WvNI/aTv0xvxWRUAM/IMBq944md6wOTdASp8ramrXQ1UvjKqPxT84qWEyfShSqqvcPEVp66IrWdk
vxn1/HR3gQbdaypRT8z4Bvrw43VttjVbhqEnSgczYIXDDrELpys54+UnWaQddrA4f6qS4KHcZD04
Mq4KO0M+jqSo/UQ49JC0cN2mFNjzQTG+jh6PdXY1MEbVYyCj+l0EJSs9ygsx8DZ/RJF7XXH45yN2
JnAj4NdBdeMcvKXF1/rK/kEL0K5N8ULfzGGFEpFf3YTGfRHLM33jFLUmqJ1d80FxJ4GrscvPgzrR
ewKf3PfrXXoQBjQ5z9QjmSPBgKiJYLzMwXJf0RDcUr+e2zWgNZ/lvAxcgKsSolccmosqCxu7i4r8
k5mR2FaMDaLC5DAJQncQz2EeWN51pMX82iQvD4gqMyR72/KOI1Yn35tSAk1359TeZ0c2l5JlTy82
nmEPjbP19uG7gKxjVtA7nK/2IBIrEYw5ytb61wSbP73X5WW3iEPg4p6BTe4W3CVU4fLNS3KJzacp
4eSuR434tjrlRjGfbVW9e5R1TS+ZmzFqgtiKREHG4e7Y/WUXxWaHOx0KsvZV7Z7+xTp9B5SFVDd2
WACLdrXU8yIJ56cOrlyxOPfzNXCCJL+TOreoCStLuLYIeTaxFnMVhgGYo4Rb1W1388nmBh8uRLOO
YKFf26IgXiffbBjiAPdXnNI316qEleva4nPG8X9pbdKMQC+wWw3us10vO6u5R9beX5z3NiZqTOW8
7n4C9sqjMWsJsGN8FTermdfJLXwaTou2lBPwdIPUrt9pQ5ba7+FadusKQMrCDvRXmfeCb2L0Nnyd
K6vwey4bABDF5R1KIX2KMmlyhCbwNJRapFE8IBEBJym3ejos8CQG1JyGI6kMswxcGkq/XWO+6+tK
6XdpJMlXtTMhI8SdF1Hs3c/cJPhso5Hj4LahQKZcIlvMw7ghxNjYYPX5oaY3UGzd3f+9jDHADMuj
tQI5Y9bBC3O187Byl1/GH3y8pPT30lwbLT0A7yJvF44/kg1hE8lJL7WzeZwgVVoDhoaQybR8wi3k
7AJglLOtq+DNDIzLeFb9RG+PVXA5CtJKdxqq3EpI9pYbycHKEkM8Z12MSN6QiSK0dzaNDXF6JCBW
fe0IbK/8Gc8dvAPYnF7kAlxAq4DMv8U1jUpMDL0kCkHTp3NIxm+epvhetHJ6UtJ/CnsynXMN+YCZ
7TRluxZgXL2dV5yGdNskU03vjOj7gwHftHSuQ+mfnpU06oU170ZkWbEZzeYAu3ZbVOzuND6iSjPs
7XKS6csXFKAheJag+AaEhuGo99GjU4450DsrvEbygcRGUMWvkQzXUoxCwUyvhuQMOnuwazmS3rvZ
S3X0N1mfsUvxtWOWyKo555vzgC6mkMfS8hQkjKXSFsVf/XPnelaIJvHVI6H9npNhBbp0zuDiFD27
6rg5hMhIJaRSBr6kKCqn4gl5gyDYPj2SgiP459EM4Q+uRYqvRd/obIbS/EsOXUbYlVzfO6GBcEMa
Tm44nMgEYAz6TnAnPSMhhEIU5CXMVanXpbABRwMtQY7rTm7VT+OooQ9kQGm/2GxdI0ILFuyZ9ft+
dsHeAex/9mw0k9upnJbjvQPtq6kxUCG887JU/noRSTLV7Vh0TjkPHvUrpP2X3UjJVYn5vOrYeL1v
Zwh5hIihd9sWuBscIKsfT2xR1+DyM1QC//lHdUL4sBQKqLA4ehReYxzRA1sl6mHzQdENHiyRjj8B
LhGk3XbJfeDy3r1uEF/S4/gL8jy4CK/1ztAfrOZc2XV3Id6up+UrY6/qiExrkP6u6Y8b2voyK13X
BjUEnAQXnwZ8mIoWW18MvkfPS9rmIZciPqy2wlEUUugQoWzoXKd9JwRn/Y/pRbEJa0q1o2TRgWd2
kRXapjE56aiQAbzZs3U3zTiNXt6nxV85CoTrkhomR2DmmMEy7I7bIoBUxFncE6WZ/hbPXgBbHYSG
h0s6Vl6YzS1SR2fH3OGL5oAGIdB+7Ao+jhYbV77tqgaoVGeqBxfmukr9t/nGG+YErpIkyTMayING
A1xZO1Sf/WjTT/SOeLKjsyHEPx5cyqYwaeeH0tis2zq7lKmQfQqZfj4dE87R22DAbEhceufq155Q
uizdID77oxBgG2e0NgJstxsgH8WXGRGP9j5pTmQ/bEtxuniFK7tFTkxhiEqlLlk7UJmaXYfKW9KD
5V/eXt7SOzSg1zW9L+9LP1/4jLpvIQ8XGyNXyWZidQv9TTyv87oqAQI3l11a6vshR3KKvQ+lJbQG
df/koXfgAkGMxf9oEacoOGuWwZ0rTkuCnn3UjZEN47oh4jddTt1pMusQ+Ky+278/vymD9/n5HbuZ
VGxKH10FYWxsW+JbePI9XygMf3sw36P1h7XV+Tjq+izUYTFsbFzWu3qA/QeMG+bydO833xAdMdVB
CtbE+LUtH82UGI/rPSyFxVqdnmkcitN09mtrOJ+TYnYxEyIgv5uWpWyfodEWqGjeMulki1t8WRFJ
uh74AsctEjB6xcKLFaQ0ov5zwjGoWmVo0Xccn9I8KzFtPyO+x8z5ciewhNfvV7HROngsfAhr0Hbp
mLnaM22Kja0lVvuFqGIAsM3Bj4mBJk778Ns/yb1hIcZNsIHX5dEQThtGvhkKPIB1Ts6ED8LTf90k
JD9z07KDQeWVtqnwUmB95ch0f3RaodYGFgGg18opzBeUBepjCaVaOYNCqCZVtoesajJfBDsuxYxP
oNDbJfC/8jnWUmgwv2WakV+N/Ipd1XvsHOkZEJXeHWOsqXo4MfTFLL1fUAe8G2pAwW+I7k/f9pEy
iYPIVbJWFCY60BedRCkMKberalNI9we5I5+Gl8NNujcW//R7meL28mfcEwetaQitaGw2W+eRxqjR
qenKl27Su8W4yeN3I63mWFDzyFB78BpdW68z5J8IjGcu86Fod6Uyx/Ezlpwpnz3ep/PLI/Byquwd
jPGm/lnaZd8bWcxCkrC64cs1BLzJSoqVTAazrJlDzH1ENeBw+HBva4JTd1wAxgk9YjoodGWlpTjo
yq2iNRQh27N0HLbMouvFvPlUbg0uqRfk3LhkkowbCLSTgQZNyQ931U6Gh45ZkyU6TM6vw4WzKQ8x
yZsFaaNdBXmHkZAMQjHOk2Eo4m0j0e7a3rDS3inuvESUD0KDx5K7v8rtXydlK5ETM4cpAmlZTz4P
GCSg97FxoVH585Y2iBossTDD+GPcLHR5WiZCwVOOvZAai6/+Jby3VWH2HLOz0OEtoNJeh07bfk6y
t43L4+MQU+Bdu8XaVb1WVrSST1+jqGzlodFIVVl9Jgt42tuz2C0lZTqeBfph5HQ3dkgkA1ocw1DE
0iuQUMfBkCqQxFWrQ9oEbzF5C2mgLIb5fKLrxVHsXJr6EFZhailFwjBqRocqQ64ueTBasD5htl+i
JkaPf6OuI21ruoDRPE0oUtXsoYoYj0Q5Gyflny45QEExVYiybY666QznBa+fnf4Ht/dtJ2uQVkWv
YYl2epHtjTEaTOVITDHawMbOvtC9tceYfRUNt2gbnZFvWXVsMyCiGzqG+U3DpWWUff11n3x5zMab
cHMBkeieUdUNb9eQG/lTzd2CcVP230lnqEmGoUGvm4C0MswHdKyuXjNpjCXYChQY8Q8bW4/5pUiX
Ga+Qw99lBSo3hKIf6EEw9WUlO+be2MymosynQvYpxesUPP35dMqM29kFfnP2fPXHU7IWcRFZv7eS
oTI6N+qAcyQWYr8BMyaH1mFk3kk1jUc4n1FOkESE4Tgo1WCdhYfMmGudcfp7741irar3x2WaUZWR
AZzjwQpcbbqyRnKkwDdZxrso9WotpprjG8ApgGTOvb+32tIi1AU/R51EsFk1a5R4+bD3KudE9ii2
dDNGDmgexdX5PBsDKt6twakQrnz0y3Z2RfjY+tN5RHMxU2ShXlmzNti1cAKFVBUHKS0SvWh8cCTZ
aBN33AgjhNyeGz/feHdfb90Py3U+5k6QOrZp+A8l2d8/crWZLPPZeTwhojoDOB4/sruIvLizkRIb
kvuCCTgpo0XdqoN3GNxECY72y7DjIsdE8Gy7xvHJq7PioaJQBmoZVFknKnYtBSb2uav4QmVCN7Ik
zQmTMND2FWaNRmZN2ZJOs9xnWm/SzNKu5l7w1RsDMIQoofm2x4K+WJxt8wL9yP+RfsIq/US/qKFq
Yvlw1ia6UHjvTsBsZoXmDYc1SJMgmPCh8P/1vNC6N2ZBjaM9M4sFbe9D68GhSq3Ge/Eo3ug+P5qx
ahE/IVv8pVeVvrEXo9IC5cNnLN87XBH8YS+BKaZCB8ITbwGLPqGEk97UwF2JxjjXUMfGNondIcSA
AeT7/eRT2VmuX8YL5LQs4XWCEQ3YFqskStMbyUrwcY6QnSVK/luZaBVX912XiwMuwOUPsrSPp1Kv
NqZW6QawrCCmYudoOdHIBz59tHjlxM2a9DW4t0tMCQIgv3Oxb5VDyu0jBm3+BrivmaGk3CEzWzMk
gwefTKb9/ScjDiKmLd1f3CWikV2+RB2BfVG2QAnhDbN2VAc5sx9NZctOlCQZj25ofs3BNyjtToEG
h/xjzSTRyOV8Xp/HoQZRyog3z68ZhxH++pKiPGeON0Wx+qpGj28Yf6Y8MaO8Wsrh6OddDLkO8ex4
Ib0i/zUT+wjPdY06hGWDgiHSMiGtmFyEPDydNYLPh9qJnSJ+vcOCrrv3YUSu7akj7Pes16E0eWIa
FWlyZfkaD74Ljh4OLNqHcMK+u70yDxR27Mu5ZoF+yveIc9Q9LOhNHiFE30jQlaBIqe5imr/Y0S8b
BXh54+C1YiAGZtAYzaFAGm/AUAKj67Sn0u+ndo0IA+3XLNLdPzxbSDQCEw5bPAGOjxWcqde1YfHq
FphlERo/qL+HCFDZ8V59htXLCsZzI+GwOorgFE2wXHeJp0a9yKsmVhxZwRLSNpA7Mrqj96i9Be5q
mTJYLNppQQSMibGMbqNqWISAfb6jh89SdgLUneAVQP1pveZz1/ObrLVrAhUETRVIcH+58DmNCrBK
P/EhQioXNqSHUC9W4kxndIbXMptndFa/B9u+HhTFUlnUAyoQKZvYTHR2hplSP9WLm25/qSEh6C4F
Wj6XtGBaVREEGqERrnKH1EXu6j0C/aBF78Jsh3QDNyNHUtX9K1sT1YSq4tPmDr+9zgQNI7cYyAXH
/vMxyEFY7N95mMAZf7V/uWvrXJ2yw7tNS5fPcgRvdVjJLGlGd9VmfF8aQyQQ1j2dZFusR3WZGHR9
VgAKuhLh3ko3qsSuXGA5iYl8nSuDI1gqyHH2um9clxip52HAY47UsaKAfgvYJw6u5HRJ3j1DW5n1
SHIym/uQbdyAOKT0RiUvATR+bfCsHYUHJYSg1CBGMx5MfD4jxngVoXKXx+HHS6o7ds+ScB3oK31w
R88xuppBBG+PbCvz9ijfWTo9pf+nNEX/AUxSABNauN43z7G3eFQz8uW/hhrnQTtljye45udkNvdc
u9J9NGEbvYIyafyEB/1nnu+luRwV3Bt0YVKf75gPFPXQJxSCAXNhG653Qrr1i+N/maeFb6Avf/XA
FV+LiY3pKspxUQWeTylRmiFgdV/zx+1RrOEFTYS954+ndu32rfHUM8nVYIgGZpAXlwpG4YwyWFt9
2/rIK9UP5HNM6MDNy9ErR8NEQ9n/mqXgeg3+vHmZkSPyohGp+oOkhck+G516XS0HctOHJ1MRqDcg
kNP9lMv/9ltMbO329ZuYHNN3TY2AZFFDRBntVXoqVaJqn44k61TLHXRLcp2eTZZgP8dRp0kUiXEN
MLnAPCbUk7R9gztI1iXfcTik7nrruTzy1mOsju22bQPNkTSrmMkslKvOSHgguqurbF8Vx+duU1Ai
Dl4UbeOoEMupfeNptoxKDelgGKtOnQ/3Sl6s1UfNceNoiF2MlG/uQGvIMF3Y+xGuBVFa0JZ2/63+
Q9CZedY/GwA6posFGig7p4pLVg2qflq4kz8mvgB/zcTK4XGENH0XghNuDoPaiC6/sTHGmnAw/2Mp
TjNQHAwvkm2Kh9qUryKKaIeB8/nn/eo9DqhRc0utr630FbQIDDsw4twXWHw3seZcynnqmFAPcfDo
WGXQPoGgJ95XCD3VOFZ38o2g2i4mfHJJaJBa68DYE9U8+kTulYCbZ5bnv0Ytd0fxQOtnSwZ04ieG
xjnc0jnl6uu26Lk37Ee8QGfrJJk8NRhLVzM+pzy89nN+0ZYNRyeuKQOzMgSxms9pOHAJ7+Vw0JTy
JQe/KMaVi1NhlMh67vbCbWFqjTPnNZTyc0LYrk++TwqTlqYrKXtXVY/S8fMDP6glhHXlT4nvkbgu
NF26zBqVZ86vgV2ZlsBaVd9HaG4ZhYo88G2GsqPdvp+YuA2e9PSWuSVoz5M51NAuvUdt2MxwLN3R
Fo6XjtJLyM61y2jCsIEvY9GxIHwlSIHqjPO/XZ0qq51IsFxja9jWF0NYXcOiwboGgA6MFbSxnXfU
3Dy4dzpq9TOM7KIMEJhZ0CaP8yN2a+PceSF0z1vIcN9sf3kfKUpahZdh6aQc4zUVgzk3Zo6QaczK
BRBosY5weyg1ZVwX85bCQ2PCJ8akjTa6qhg1LCUm6UqosX73QPqDNfAjAi+td2W8auAYFWZ3bDRl
XHr7g/LXGUGZ2EDkr+EK2gyMwMxGMWBZCoDqYVU3VaZXqct9UeETdfRQsZkZThNTGpTqtLim0703
REP7H+gLiE/ZkWL/XMZ6LwEJ045b9eXMbhptbbjuyMI6/QUhXjwAOOTzRW7XxuJ59wyTDYsgphWk
oMo3qSpkjoGShJL0gq0HoBwEc7TBYj+XsEYxPggVJF1cw9dF2FbEKa6HOOcSN7v7JLT8E70CE73O
z3zVpq/QeNjALPQQt9NoukV9p++HfeYkjOq5nF9sbL1EvV2EN16GVWB+KC/Jd2irwsfUshvIMSJ3
Kl1GKmLGZxv+NijlTDzjxJYyXeGbkwfjW3Uk/89+tuIGCVOaI0zHFKPUzun0b55RpQjbDVVWlXR3
l9Z3JC2DPEHuziczEfGFI/tZ9RgZaDZ1LtDC4hOojh71VqhW5/WOqBA3u8d4L4hq9egn40Yo6exV
oyVQKydzP9u5eGoIfaPiUBdcBD/E2zW2rduaY9A7w8TSs99LsuWJ20G811pdsm3w7Yu+qwHa/P9n
6G90aBjoFMpA5ezYbv2bct554dUShtHFsaw1EdnsJ8opHHBoMWL7tndUqJ59vQyH72FbQpgeQW11
dydX6BYp1phangnWDGnATVr68cSdr/hzd/7jn5CBT1Xu6Msvg3rL9PympClUErldPU/6VH/IR1vB
PnK+beTPvwKygVhE0Jq8sLC4DhzgPrUY31eEYge+LlWym+ex8xPN6ZZ4NX/jqrW9WFF4Vp7seHoU
yLbjwlc/l8Y1cdCnkv8MyAzG+IMGZE8ht9J1JxebUgDyIg9lWnFc7n5e8NJ55wX+G9AnoMLNOcsf
L3jDIneN+kiiQoH9784krBzUk+m39LiVOICWpImM1W/6c05c4hSrizLiAGze24p74XD0t/Mz9zcZ
fhGbOgdraOM2ct4lGGrSzN0Humggg3qrS2lDy3rnJFd+EwT8LchVOLOVRmbgRib2YEslVp4PjXce
8VrdTcuDrDlMrPnlNBpTdqpMFkqSXEUZ2QpQx8wNA0hJWbJ/7zrq3KW2bRYLmC+Qb7jRxEsTxwdb
eonSTCJadNWIk5Wnj+OWtvV1lsOYZgCR90iSgEjwjiyr01+uODC9/ecEc2qEu6fUhFvq/NlBV3Av
cN39206kqPO10sv8qFAVlhgsH7rAegjiRVx5RKBtnkeadKSJ8Tm52oDDzhb5XW2MKf03NBtZU0Fs
qMpUfwRcZeprV6VEsgZ787E1ocbPTsZLCTjvVpvOKAQRqhLHBaoVwWHnyZkQ4OxlPXExbF7IJHi7
w2lWiX363z853hbTLrKUksepG7T8/iS8X2ZNiGLjT+Yt86YieaBrblwW9FUUhR5PQcFOw6kAJRgB
vVQCfBkl0AZg/2eo/gd+vVV7fqoNbkla+4ADLYAc01baZ6KxzQcUplFe3qppBZNdw7ZX5Bu0zuLT
TzzsBlwgo1xMnJ7ALvBkzOry5ugy5s+Qctg34l6S+1KgQB6DAf7ZwEcamHaYpUBLzgNAq8zKcLQE
WbIZK/DTyVvQ/3K6nf9Iy68ORjMFcslir2MYmbQ60f81SWZlHUY7WmeKe+r095DDIffZ6zq9DN+e
CSnnj7AgU6hg4k11LljQMc8j5zlzx1g/N6/m7i8TjuMTnHQCWYCQ1Zw4ibCsxBvpmVmp1HTOJQdn
AuK1uy91aT6OslddQ8OTUhqEl7TOJ37n3heFOrzNnstUrbVDjLMBEYuEtx0iZRqsrBl8+Q9GZlP1
M4F2a2PQVUxxcqJl81ROp4wWxL991bqQTIpxtAIoiVeqJtVBdrCimcdxOE/666gABnYYvcFpCBqF
sHGHZP9Umcb3YQnMz4XlEkuTiGIurRreCuI8lyfUXSnmRv7U6xtL7DZONYXGA6xACovwTGFvm69w
Imi+nENq8ThYm6CmQZFHaBv2Uy8cCUw/PfstMvfDJeZdVDrJuCIdlnKakKWvjnKwdALmJJyEuVHF
VdNASVph7hdAMmq+GczOiU8IPHnvUhRpcjKDuSjgyrHiDkCQtFwqrDAOyWXBfmROCIJ+qUwHh1iU
+20mWZ1vueB47yuWtD4N7RU+KzHerKEHZANp9K5eTrstyI3EDkc/GP9ENLeEsGBY5jIn4YbI62y8
VI6aCyLPtNUVzeLP5yCzRQcBBalVFmB4u5h+8dbf6T+DP6mOM0cN+snNvdJiWx6EypuLyQIPJxbf
9LOia3+S4Jgpl3txN3A151ipQbyLR5q/cC0YgmxH+16ys6ncT9gP3KUnEbleadO71hKZZVfqQagl
PMOhjpeUdJJ6yyrM/OculyS+EMgYzo6ETPu8HHwW6P6obA0on/qkmk6HqGm6DvQaZ+/6TPbUk78C
5MSXOjSM3gOvJ6euGpYoMmQvES9q0a7uUY1NTVko95nhm9dgOx+wo1FzNUQcaHOn+U3lLGj6pns/
rPZLP6EudGy9hVHucxJGY3WLE5leUdlzU7f4NdcD0ydkJD4sMT+hVT3UhgMS4K6uVsqy3ClNra8m
unHkGUr7V5843JizLGfOnAGS6wL1UMFh32h70mYavMss/pP/LREZBsOrt5R2TWb39h6k8ACL3A2y
aukr1NQPa9FzgDTqDVisRl2ktZNAHVkMk9nBPpv4yZJssM7yJQuQVoWOszv5FlyA5gAbat0k+4p7
n4DiFR9a2+3t/Wv/E6JsOZcLi2HJeCnRhKJ2OK7LlB9SULGYnUaFYixQb2MUh4ihtTkkdDiZ9Tms
8x3Vb7Moh6p817El+0Iv744Tp5amdK5IsOJ+e/bWP0nil0R9MoC/7EFb2ohCh2j43haJ65x/HSXW
Pp48xCGa1UHQpYewBNjN1gd2GC5Cz8kyzL61P1dpDTkoe56MqbjxAAEMELPEQKx7OIevtoIr0fiS
Iun2FwtohvDoE44qJ8Hjqy6RExNM7IA+5fMShegTl2vNuApckyMirSSNgz4zAEtmOsY4Od3lLLmC
8MTqW1odueAAVv13ygEHYjqOeqtsee/w/VdEQoxYHfCbhT44S2XC8lsuPMvSYfvTPLrCwiTo8htK
rgBOMvnRRu1IfWGSO5946VH87IQ3oUzzpcH//Y1K3fN7LzcPyR7v5z4QSTERFJzUnZjNVYl9nBuX
Edp0SauTdSbGGzPHVhqSdTId2RQI28r5c7QuhZ5q36LxtnKdM07a7kpuaJHTcjN0cTZuTMxGZ8ri
0zqge4+BHbSVcERzRKysA09H7Ki4Chvn8bzgfKPD7tE8ijws4086Paw4JX77oZ6Tb5vBcKNYYHTu
s9VXSwCKysBfcX7eXga3NUW1f3fN0VE1Ufv4YI+FqB0La1OZHUHrs3halifzE8x2NXJFPrkiv3Pi
FfN9sjD3cLXK8dOmGCl6vXep8nDtnCMzbQxY7v+HGhxJyJgZhuCPfK+kyLVD49oKA3JsV6xTDWKn
EudXB+kxt6HgS3lJmMH+H6MWYpllukOqz82bMwDCByXGXIrS3004GV52GWPwpDgM2jsac5mepfHY
1qcqHeTf3RFGVKZt4qfBHSwvsXxCwU0hh9xJreAPVCOSih1PRMtTZ0Mw6XODvSzhIDHWgt/1UvP+
vP+SrrnZhgrz+5QSf54NxjshNIsb5ztGqqu36iw+7IMp3MEhP+XuzbOGuvqWTKnXE/BAZ3jn0KYL
FkBCzvsb7h0VaI8YnYb9ytPk+gf/CwmBPSD6bWGlNi/46IWST9v3UgF3GynT/PMe02NN8FOXMZq+
hiKVi0vhErpr6bGrndEvfODJDOC/LIiju5jVY5h/pIfziy6YqWYw/EduI4Awjij2CG8SjpGj/xZC
+4PQd9wvhO9M/JvuZwdRY9LwJLRsu4XuWllgQUIVo4QxPJSCrj5bxq/YoppvC6PhV/oYcTS2MVXZ
zHcuIxbS4ohulcggEuFMFpDlskTgd6Y8rahWiZzwnWTfS927Zs4abTNwBhxfIuTvhgdqe7lJCc7u
FI/tP7aI8ZxbnNG18EkITWkxGWyO5ew1BXHbqlD9+i08G7kGPlNKpIrE5cS0CcCV1n3CmYaBjT1F
B+F+ud3k05z88IZ46FowgtiNd0CrqMKBC3x+nHi2Z9Xq3vRU5QuIVacqL5GJy1OUtT3TV1vBt2jn
6t+oaxx9tO9T5kzEIOH4AmksIgAoHyLjQrhbZO5NGFxSQ/L6PXUaX23ku9OopvWyPve3xlg9zq3Y
QdYKQpCMAfMofKhHzM36LpT9dz8V9bO4TYmJdQRpN3IpuXhtBq0+jmQfoBanrnoLIMtwAlHB8xpc
Bb+bU25WKJijcKdSLl3G9AXr2fsplejOGmzE3qsXgGzlcvJGuWrsK7xpD5eFonvG1r0O9kK1gqxi
TB7JMLHkCkKLqtDisWCXn5iWPJFbCIB0zagnHa48vv7uWYwDAfJZmAcJPaOjdNN+LaGzySzq3q1u
MY/iocyUcXDWz/hnU8I0ymCJH+AxTHEVUbydvczJQUFNPKUVs0+7obnMY7CCuSeg8d26ktpchkfm
8mcLmlViIEy9Wxg5TX0vEvh5DhoKuXUWB7iq4cstZsCt4QkzY1nIbppWWemyuwmbcctOkqYM1nE1
E/38pgO1zHgbXdOP+GvYmR4EM/eBH6xEZx9AZ89oPeYbvpjuC81f/gDiruf2Xfm3uMZjAQxm/UjT
2rBm76hn+G3WBiJIQagL8NwIq0f9Ne+VFXsEGlR2SSc71q+Mb8KP9QG9mfd8s/DdesegK+xzz5Ue
4TnjuXhq9om2kJMypGjdOdxZW1t/5iEMgmjjvD15/2GjCy8WzjKBNyQ4qEAkDUFlRjFFRvM8A++C
jKKofVMZgmdycepkoIBwhg3sCwGnWS/UrOgnxBW7yVs8rpFT1npaSTEk+nP3RXJ3V0Arv51IPYVd
IYKmYy/qx8Z7ufEMqMO/mrd1jBx4fW8SdTn6PRzbPVO3tXk6nFi9VO1Qj9pyhcItEHqlxiibiq3F
F32Vuu65EpAZSS+4zSA8sG7vZqvr+vvdyfO3+AIkmbfv4+4YTuBWdrZfqN9WFyN5fweLjYiIGsJd
/I+X6OteC6tUk8xLg9UAfXxkaAhwU+h9MFKFjFWIY/+Ntr5j6D4gxa629AbKVgJuUDcVbmZJYOdC
xyslrmrpQchSkb2k+l+lnl8X1zcIZ4Cr5nPwMmMvb3TzgevGPKKqmHbQNqubuqQjJfg5I4+8DHFS
MoDVon1x5OUyrv9husUtcpWY9AB7hG2x3ZqW1/nwLn6L3A8rVv9ScrbJG0LNZHp3Q8ma45pX0m/X
B+uJQLPx6mdwnDnta6adZdav437vFKYiWUcpUJeECEilMcKz3qQAMD+CMD3FSc2ezarTWcfypFFa
J0hS1X7ma/swji65wvryUNPThWSqPQohS2uyTh9sMOYtihhy2wPbTBVUeD1VHPfkqvK5/xFjOZGb
IxrLovgx9Xc2GbgZUNf/MwptfHheN7OqsuZpObtZjaSgZ3QP1WWmUIMIFf6dRn2B2tTqKKGJWbcm
nAUNqUMAUUf8tmpgtD/Au63ipE0YUqNAFyVDvogy0v7oxo3UsBrtxhMdQqwqdySiLo/GfbC+eeMk
hoTCWSotcfaM07Yh28th+ui4tLI4kOk2QT1F6Q+Y3GUusmQf51FdYpiShc+K2Yf1JK6/r+s4yzxw
JagJpnagTAtfgheAPdMwMhuGMOI/n45dTpSiyb8S/GOiTg9MwIdvjpQAklCTBsQnaNNTan04WhNw
Yy9Q+JX5RA/lCBxVNvYXJoU3CvY9b3IFmUDFw/0pqdKNwMDIPyRkGRTpiXG/wsVJ8HbaBxN7KP1W
YWv0TKsy2qQMxNXnC6tkJkM/Ss4Wta2QsZWN6hLDb93H3bwU6P2/96KgxV5V2snULimoovA6eXxE
u9q7uuR4PNxY7eZTFvrpWyYzd8QPh7XjTwHMTXYEiEeif6NwOzp5lbP0Wgc6xEoYvCKGljkzklr/
e4nbql3hamhCU1c7wx0eWiQ5sGQ60NMYo+U4pJdHrX3aD3OTOR7HIaOx9FiW6wNQtl0HH7TOXYzb
3jz0UMfAsdumMVwaSuGpLs0HDL5yYezsjBpFaXR5+uDR2q2GsVO0bxeEympdELWlc8IqalmH9k2W
I1zxHEHxaUf2g4E7leYCQ7E+shCpCKRdPuKytbo+f6NZ8yCf0XLyLvDh2ZQ0edv80IZ8Iq90Ff4t
vJY9Ln8ptHd+58BfqBxDdDN6VhnrdV/OQ/tM/Rbc2+uSMmwXtxZq7j9fBK/JOZm98SjVDiK5rmuw
1EVG6JLgXDvBMMzxxmduDdbPLdXQhz/Rlgi9ME7B5nnV1b4Pw7tC8fNM6B49POEumZNdZSGuIOye
9+jJoMZEKAYa6uffbIRwdX2nhZendw5Cl0SpSayPk0yX2S8eaN6V4C0ZgTFcMREdr3fYvoebtRSX
C5F1F2lLqtuxpJVzcc1sWhJPZmdkTm8VaCM3plj7HeWf/TH0FeOzVc1LbvDcQzRoTu1R8xjxag/U
kDj9QZK94DwtD9if176h0s1dmhjA/md+rIJu6AqUMjbYRhRXTBrSBVYepSa7EfZZ8QlvsgXVUto1
Bj1bZm/TsCqFC0Fbmi8kCRS19kjF9DQGT1N84BNNR4EBE9RnKmDOA0FKupRmsGt+vsVS2LZ4wuQI
Hyg84QHs8wnS2jT4JWFvuNmgPAuoeIqMtGwAtye0gwJFfPv8uEPwZLKRFSfCaNanXMuYefbvmou3
C9qsEGk1/OJYXVBajNUglcjeM7Xl6DRuXVXdCLWfbdsSjFI6gJ4oNhifheMCZx5MlzdKT6fX7Scq
JTCQ7P5MCwaiDQbtBJauiUt4+FUez6rmZDyEKp9RviL6DGtTeSzhi6J2rCMvDrQHdI62cnogFCIw
ShjYJDGv2cYKzwGXQhcu6E2OFdekkLtf2Dqg5qqYtkwoDSBGPLd0ARe1QflMF976bwhh+6tclj3w
NJZAYErUKCIG8gfdyAXZvu/Lde6AymXtGEEDcwxM6KN4wdCJ3VXbRV38Qdsnk9vscpxlxyBuAXRT
8XkGrbJtLCTzLjNZoKbtrYUPIemt3M7WjqvYpNcOcKocpPn3S2r7MdLfl+pF1RSuK9jt8C3Bkm8Y
u7rsXHKcy5ZlfOdsRfCekHjzViQPawqawwnLA1q9SkaFRwku6bI0tNKsgqb3MA/RDonl8n/TpFOF
mWw2TbQKv6t7oV7PxPTNTn3wa78dMGJBt6JgNreneNbWd125vgIrLsTaHr/QSs3PSENB2oy4uqzV
f+nyeJgq97dvBoQDO1zcjiux2fxx4tTqCG3CQ3/tOGocanB0u3fGLjoIPYzVxQUmiGJGEvHRsXdy
3pkp30fkBJwT5JXlWqwFykxVkLj7K+fpTwwJifnsVL4EJxEOq/HOvDQF5uxwiC/qGuVKTEF3UNFt
khx+wVDX9GnSPyEwIMUB6nu07mbSpbRDukJywtn2AASVPPmeDT6iQLD3C/CZznlyjdMb39hNFgiI
CfD+XRMCvxJhSdVCPErX0/Vc3btMJTtUY9dqRagU98HzrhHtB839Y5NuxWFLauAqXMkmdxPDuSmv
SzNChc8Orrcwy7DPa9SrE8FwCx9e8a1/x4TgzgPC4Qv0QFpyJogLdoqh8bvvAffYaZCI0uZIlNIN
xSELEhUdCqz+4r6bvGTgmMjuHnxy70/oADN1m2Lx7qDB1b+Bzea1W4ziW5kYY9O1/XW3bUtVWRNR
CO/p9Xcul/+veeMlmO8xl2AlDLt6wmLxX83MgOXSUn30Ls428tsyUmjN0Y85vDNJdxBluAfZQBoM
dKRQS4ywVR/oMDOy/F613+NkGxbuQfUpfqoYXP7mtLgeJxc3GEjvtBe/2p1E7RpUqfoW6v8KGMjT
/Xm1ulxFX0iqmGX7RkyR4tczmbX+/FSlUe5a29s4QhTf7iNC/Blf7kL80m/Zrt83qZv+If97MI2o
i1IK1rf+F7yRyxvL/2LF/eyOciU8h/XmqrrOHQ9jb6wxm0JXXieRsTumNKG9rNWj+aEKkE+9cl3c
vmw9PtQNvPv/yOeYyfaHnAwZoxp8/ok3+ARwTJGi2YDWtek4Xrqk35+14oqrw95gbW3XvqdU+XkN
zbP2B0huTHpXDXLJeHQgkI/JZhYRz89u4cKgM3Ory/oJjDfo5R8SEuEQNOBFQeDFIjXICM0HfBLC
h2z4WMopcXosfABH4zLOcpw/KklnvONXjtPshZb2xtGwBcI2wL1K6LBVm1J3DlSb0m+yiRCOTyhs
Xp9ZQRJ2aMH6tdKLhAiA4VLX7DqNHr45yxxIV9uAr5zKnWLD15LdmCOJlGHxHaVaLEoZgKxZaOeQ
bPTR0fZHWsvI3+Ldkqaj/rVmMgoHBl9dgMrWUfwprRVH8GmUKgBj+ERPFSURET+ixwOjN7Cmy9/Q
T3mkzC5dKRdZW1+iH5k+LilmJl3dxYl6xUjuw9Hkj6yQu4RXKqIiM5mWK2JGlxTSN/3PvWGRmMgM
4zgC9dOArLyF/0Q8N3/LoERW3wJEUOQ516kIW2WsXx3EDi3GFMxpAqbdi2UOiSvNpfgj2dpOMPPq
TiBG3GK8B7eaydGUA/mHdM2+nqqgx/bcL3IUE6U3OktB3q1E2dWRB2ES0fCYQUgXNBqDY+LwInLZ
X3VTx6E0rW89G9OD9sDrokh4iiZczYGVeXL4SkILNcNshePCs8iDenScBRwwQbbusPnlF96Mc9UP
p1L3aWFeOJfy2yak/lk7Y2ZpavWfyVwrMTUxMXSlHyubZ0DbLYNI7ygfTPvpNiKxhALQ+BXQwgGw
M6aOU+ssbMGU370JgCWO99+G9qjaAmVP0blryJzDXzjqLg+vsLLnz0aBVkWTYfGLtH2jiNuXU+Qd
u4YsbZuTl/89BVX9eAMMXVK3c6Yfe2EXHoU9JIivyCOTwVX826XU2bIM+cNUyQX91SOQQY8WOj3V
IuFlnCBOXBIll4jlOKo1nEW++Pko/BW8qFq4RglOHdfOItTvOUYUl+q0IHsZ7PPX9Ecfpm0KDDxI
9m3M3UJ2Zeb5Q24DuyJxex+ErFA/MGOModkc7gZC1/mQjIRe86JQH5ylz8B5s8rduLcD9iadVEWv
H4DJ2u6hg+SDMgjA1zf/kuUAPjG+5h8xOcq6Fsgr2Yvoc4Um8hrq92mNutsAuadtVULp/ezpBVCJ
zy/wipOg9w99d/cb/3RNOWRSAysAJp0tAVJEvwlTpfso6RT2atujSIGGQ7/oUqWenJr/alTK2r/X
wlLua/ZIgmI1v2wXG3w0LcJ+zNjZRDwQXzIPQa7Nlwm5sRwlSrTGMphqlJFNXpD6Qx9N9fwfYddV
3W2gcFn5IW+dVVxzOpg7mYpL6k0CuvEaNoOdYjofXFMU7ykMVEFJDBNEYZJTZBtTlKB4BN6OlUua
eBETNGmgdpxB4agVH5fHwljIUR18GmxsCy02eIdoi6VbWOb7AJCc+evQ960NJSIjADcRxP5y30kP
18XeFj9OJNjh9/JCtWpqL44Jyde0v+HrThjzIQbrkwKqQKJpSvOj6HLC7FSiaGd+xCwxovpjfHMY
htE6lQZSlUn+jQz15RYUvWJkfGQblMoY+k/dVaKSaiSG86P32Jv8rUv0QSOxdQdxLCHmf9NBzvjm
V/weGnfnbsphjUAKel5+cz9qvRDs5yvumcs8DuRWHfDVi9P/2Gx/tMnmYrw5a8wFJmcAZliX1L7z
ahL39NzhnpGudE6zdnYq/nv97QI79kAfyV3jmzw2in4I8Q2OwXGw2ybEOMTHjMyDWub9RbSeetNd
MJk+jTVBShU4Oe205r6ngUyCYsacaNdmmT2PtTfGrasG/kBJL6yXlT9FCqbSoB6YQcns3hzPL2pL
4XloMVoBjBJRivDzdeNnQFW2zEQj0eO5VZTKHY+BNz1NyzQ9fmuDBgP0GBmctHaMU9BR901mg4dq
JClzCTBiuLSWehKIGGDqiz1/Ft4VS/E5J2EpXZRwMU5YBl82LksuKybMUCNOSoOJi/JY/vg6xUlm
YecIxHApkOdHeyGleWwgxnMNQNG+bj/QBCNGoZUlpDAm490hQOX0sktLlJttRlORKVy02AbGjkfk
hni8VlqL9DldtqXnTMUgInJbm+QcTaLA2uHVcTPO4KHL8ygsZB69N9pxx0u5zSLolKFG6psceeCI
kF00uL8wwDpR9kkJtRWQy2nOmgtm0T8d6kxOrdKIx77lf+z6P8SWppTXJ8NtyW9/2UevfO6U5t89
BkbCdmfmKVzKebqiQMUsRkG9cQ/+EDw4UTro4PdkD8cQBiV2XvM/JpwQ5IMs8IYL/mU/zQzM+Olh
vZI5CrcwgTqUUM1PSoaNcxxNjfqPfgpckbTPcp9oz2b5ZrpMKyo8grlZ/GpnD148Dq7Vo2GVl+qg
MvnM7x0Y3i8nHXBXXylJiw2yksNFrdZ1EmSYaneruxBvfanW80a3KZqzApWKJU8PCZn0n7/P62lF
jZ+0y0sL3JKSc4kfMpXYOtVN+UIFnQ9Tj7CRvKjqJkavQrhfteKWpsU61qQOt6hfZSKrvAO0c5ck
MPykyHbCf4kKKyMwfFNVFqHWj3ge1xxJ92PBI5KYtxjBfCwhSe7eFoXeug6zYiZWMSLNH7T8NrvR
t8jlZlx2GkXpMPksYF0h5hICT4tPvBOHMqLXmw5pDrvhTRl2BgoFND0yc65jaJIT4IOgoLWlQnzJ
jnE4Z9Uwtccas6xwQOzxdafZjMqjZi6Pz8GXNedipROjj3ASZUuh3vfNkob2R0KMqkow77ICzR1N
ETDXprmnXkXMZ3HjUSFpPpsAB9lpZ3FUhpKodVKcNS0PvETyZqeD0J3T579orQNRx84cWTW6NG57
6mC2bH0dLu6PwOgRKxrgRt8CIoyhNlVhm9xp4+bpww90uOtXF5pZtIFvUH+rguXU+/P25pjlU5Is
Yl+e06dA6KRnVjXVjPYSNmfG1qx7FeO2n0xuzlj2KgQ4KYDFLLBx8DW5TVkABBhcONa4iZ64DNvu
QD1q8e/v+sZ5eAuc9sHsbGPZDhS9npRidSSCAULcS5fPpQG9TZBAMI+DFGTrpZHZx/4ZUQ0NWVde
vSR8DtMIkrar3PJeUuSMhHgykL8yiXDzZ4M/8/4hRiywqzJRDkSlecGVrjtu0yjLsCTvuc7xKM75
g1qQ85m6MBGmzt8N/5kgXg5mYHPGVHA3yNTWyUNXSni3tQq0DFfJIbZMM138EX1vmzFJ6uj3y0H+
ZzAbFqRTrqLZdWd6j59UtnzmYCHGe8jPVGVL3jab2ThR3yP85+f2oSbyZfV4sonvca+ZOlpEuEfC
no6jSD0I+bIofdER5O4ZoU2P7fqf8I8yrG6GG8dQlw7/1fD6NLLw1mAjLWsWz9+s7C55MTn+BNsQ
tB4cxY9BPbSplTGhLh4Lcdyux1hRl71G5jHbF2PMOhaRhN+RuNFwE6nV/cJHShN/GnDmYZIdUNsC
f6u3cNBTBF/ExO0b1u3RUxeTa+ORmcB5E0YOPd6MYaBcqAaSJZ3hIKEfnBsQJiB8GIeHGtVEmNMd
7SeqzObs5bztzwpK2GwWcdrDcpNQ0NoyPqsF2h6T5Covz84a7PwxN2Vt/vzZE5kuPuGjUbxsNjbH
tL2Q8/e52EODycTC+liTo39jfKUc3Jf/StRxq8PsMbUHBuCvSmG5VRac/BaQQot4XEf75+9h6tEA
wfAEafQKxMcyrJhToxAsJSPdJYbATbd1lI4y8TxZVVinRmA69/deF/nPzkm0xkvxwAQMi7pqmYjm
dBimd/JpGv2+kP4QzdgPidp5nEhx4vWPlNNnQ2WCAK1sYc5BpJgBSAlJsXluDg78rR8rbiEp9ioy
jdJGMpiqNTiXEVHCUbyuzuVhq7Y4KhzSEIZ5ADGQpwBVtoG+E7cszjvQWp+GdESxNlm6E9ouEfYE
Iiguxlz3CfyshD6v+mk/hLRY1uMVulFTMPgItUHOkKl7dmmYJs3tud5as1x/VN65CKlENDkegkQf
hfGrJqKl+u6+bSu6NriIe4w62nlF0rCvAHWpNU9H+CxTJp07WUMMQcOfL6QIsZm/S0oEB5hZnRzq
naFY2RnC7E5xJmb1z0rclvciCYcAAmTKJjDjO9N9bF08Cjddqwvvv99F+kHzrZV0nZKuUZ5GP+ic
/v4IpTMxKtESZCzAtwxnhLfaG/tcKahcLw3W06FZ8xANUSqcnt3PK2akpZAPiLnlrGNNH/Cn4g3k
YiJ3VfZixshN/nWQCJoJ3eY8VPj2Y6EUUgPcBYfKdJHRXqRfk/gA4gl4J/hQZHaCqF8R3Ep3AW5T
s5v0Fyr6WspsVeuNrWpps8szhBJhpE+1eEnLW/w3rZpJYicGuubtpwCg6rmSPwM3i2CYItKNkBZ2
Xc4j4Y5CJDRwAMBf4ybxNvrjJhfvss44ojtqDiacO/4aNJDVb8qKBd+FPJ/fREP/XWzv1soTlaVm
cNIIUCmhYYL/JgS4LTE03QeIkRgfbn8ifFtJBpbIJk3QCtXvolPHazJa168Urf+BD2rOOZH60FJ1
6MTd8pc6CvOO8rOyixBT3k6EYgzzlDk370zJeG9ahlkd3sZV7yAPLkFr35it7JnZir7pRcKjE8mY
vPt2tTo5c9t0TCd2Zhpxb21VfZxCBMH6U6LBOwdWdPMXARN1eMmod2P+GL/cX3q+J/o5dnGaRVsl
S0nxa36QLXN447hsBb8NdvUELJWXhaBNQ+0mk725mmmMRiM5WKBMRRm1NjL3Lglz8d5/NG5OuOsW
mZBPhBECSMiHgdSceMp/ilpgVuYYptpOmDb7vsJbQ/tzWQsVJvigZJehtH2UXbT39DAy4CjU7Grv
3cflRdjjsMBmfSDFpJJf/g7a+x/+MEdri4ziG3j8XAsirWwM5jbMwAKoqZXmqZ8LyS9OZAxE+W/c
0qH85/cMMfHJgSCh6X7pEqTioclj+tHNt2/mmtnrBLvhTNpCmrA39EyjbYm/V33hdT+SM2t8b9aW
bJ6ITpg7Wt+UMmxgptvU2cc3q4VQDnNBrJ3HXpA71PZJaE/5U0cO6xkRun8mw4SbW+JFikQxgFsT
06DB1L3iQFBj2J3AIsBNcmuU6S3liHWFFtWuOkEKTJNOnQn9WnFqSe2oSCtE8+CqO5MYufI8jNk5
LjlRsnTFRGd7c7g2CFO4r+7Scbmck4PfdffYyBtbA0MXnAoanYyvsMaPD9a2k0Vcsm8rozpTULe+
VD/km/CE7CD3z36j14Ab5WQF/k/Oj0I25SapUrQRhAo2aZjhK+e8HLMDoj1yzoCAfKzNoCdlaSsI
76HBVXs89SYs73Na3UJnbnvGsXzQhvgUzmwhDllNUy2zfWjNddgqki/b/Tno6nGjfwFYT2rxBacI
/hrlHvERLibyjTyUGDjKnTCKEzKZo0KOrRQJB7tMnMkmk2Hi1csWOIikPq2U7G/yBUS/PRtHA+A+
FH2VF7z6+bB64KnVFwiOGFxv1EtH+IfIAOKvhDb1FAxHyKigqs3ycKprRjIwIFfQdDrZiYKtdCDR
S//3424BHqzAdMsr0wqZuoZPsBD+EI1wCVGI/JPh8H7gYZCMtatXYTsksFjAt6N1iBYL6tdUqbFk
M9ERNmrrepKrZ3FabFIieZtdEVeh5F4nicIKkCoyxNZ3YkEZ+bCpITs1MxtEOqwvyhfXy/vYse9n
Oh6hjUX23zSufsrCZhW6FvgbMKzPZppP/rMzM4DdtjRvFZcQetis1YCltHeXkO1+h3Nl35dsbOE/
567WMvAPB4foJorMRz908U8X/E46O40EZuZNAjaeDsOWp3+znRiAlMcW7RDzaLgjDqI9rrLMpve6
JoEc+rOaujcsFuG8itgnym760gEgL6Y8oC2NEXHKQF7Uj5xNuxj2v8qzud+HR85El0tQrB3EjM0G
XWqeppa/i3bUI/LouN0tWSDgrFNWr0rVH2vbuBZ+Q/5uwFR3+88Gv1uymhOQAKhiF6JRSMPn+73N
EmCN5INsJb/3rOjCgy3plK4D+iYoIzFSIIpc/+5rDwJGocXCXnYzOWjKuDzOKMSxH2BnyT+ya08q
99rgSeWqI4zsvkksUe/DawCQ1yTmePMXYHq5GQSgPxvYUp/hCjuYRXcnr0X+Z/N8r4d9f/Ifewnb
9y+WqDjYbcygIEHToN6hvhFkLqo8RAzji5Tzt7W18v633qF7i3PYVLEqaQqTSb9iO6gNMVVycEF6
YepXeFFq94v695U1hojeRznKflwBCoKIC9Dse47XwSctDiaJjW5oIvMdrDsFNHlmCTHx+WEds8+E
iT255PexNJTc1MTs0GUPEnxwBeb+DQ5w+rzu5DRBAmNQsnhnNvDZouDk/4ehCaCpmVUoEIgfPQsT
58ZEC1+pgb8CNderZdi22xRXP9R4Wtvh4jkE/68e1omdsg+GzGlubxqP+sYMsg5MxlEdh3xzzAMK
00vGyc9G1C7VXk6UmFg6HuXWrl+1ZUa5z/kt88RFP9rbFSK1EJCgKpS4gq+lM+B4YPEGw877UWqE
OUvO5rnxzXLEUjuNmV9kAqEIa6AjrdPNHMpvyQlaqqp+jvjyZvPAW0zLAUxcHCv5S2yb2GoyFwgq
MAXDlWOJDYqPs6Zsd/lBXpsmaBJiIIE6NRiYbIY6FI3xjP8CkXGyOwfNwDhGTIvE1fJd76qJlE8F
EkDOGYhQ2m3b13R3sww0ywuiIjwlRPT8bBlPVMAn36Ur2whrckUD915bnHtE37/NZjtYY/D2HhwL
1c3iKsg9gx7CGKeIX3RdX4tyEroqdxfwo/8biNT6KQ6HTj4j5g+1k4AQxofK09o2++k7sc6JU08K
38Kt6QobEafSv1D7aM0H5ueiZS0sX7gwPwjqlxKwi6ULyLcC90F7pZ35viDbCTUPSM8tHt8l9A5w
GcfAy96l2YLXyn/5J/d/esK5QsnXJhLq3k51ynESu/zVAiMy8sz7TnkwUScjHpV0iir3+iJyeLfY
p+fUkXaJRiFe/UT3ijs1cmF90TrtRLFRKpctCxxauPoeWdDxUQFAIH7dBMeuWcBnf3sL751q9WY3
0VkCG7yL10lI26MSklYiQPwINEiOJn9ZMLZg+pN2e1r0nMaVsTCh38pIVDCo2fwlmKioplml2JS9
rJBeRNSUB+XB0axIdk/nFvKvuXfrEr5AMc1tOADinEI+Adz7j6W3+C3mMYi6YQ4gaRysOsvXVh8r
SpnCyqsccc7jmhkBmN48j80ZCZH8T8up2KEgrJBriSrj0OAgTwHtaPNOREzKFCO3N6EAZvxXgWPk
ThL5tM4FjMyGac2n6048xG1vLKZlP3dxll7yLmPvAnOWyAPIUBhs160mCZ2cEJKpLwK6q5AGZMPS
Pzahz/ne+8onuNVpKUx8iEXe128X312yd92ciyl1lCMbd29QAkQg4L8jZJ3p13kPNILQZCChQ4zB
+ykhq1PFTbG1OqV/Z3poPm0w2EnhIbQ4Q9B7ccGCIgOgbxjZtC2LJR/Af26rdt+Z++pcGJsQwuXc
zFCzVeHuHPAIBki8xXFI06Z/g9PgekAdC4WR/8xfOtdRrX2tYFZkz0DTdGZOmTNitY+HGniYQXIY
DoQrjwwxuygzMCemJiK9qPoDAiDO6xF2zmuSxvD/2/CeaeIsQjpZAnLSvzjTK0oo+/j5ySwcdSeR
i4SN54JJWDiShmDtCMtVRTquAk9Rk8qbPbdlNnFkWLn7CBcZOrsGpNrUwX2NNiHUAabnESdyfkvi
bOT8nd6CzOlxsQKgeSxwQkKPjlE82rfHm7RCjRON3niMSuoobfe2pNAAZ6L2X6nAkGx0t0KjcStz
5Key/EXj1b6N+zJ6aksh9aUtbPZlK+9dDLzY+tl80Rf9pptPGRC2WqbpXHvH3vFLkPynttkdkmJs
L4fRbO6597VE64QabikAatRru537cqkt+l6spAZVJRUj8UnQoRmHysPVSQDVXvysm23IBUkNYfgG
PnIBKyhct5VIxKHgIyRLxpD9K++3DlUpDrH9VOPQ3zSAnxpiY0x/pHmSC9+l9KEJX2aR0oPuJ/J0
07Xu92itBo7ypCw880iCBKOXfRC1sHbhaPqLiXMMzqXDfAvoYI3dilhTX25wWSEJlfArdApVXLj8
K0+n22aHeytSRCaivwaqiuZHgHQhD/x3CyTEju2KA9e13quUUZGFLITORqocMAsIAlcG7YLfbMGG
wk0Eaki5YUoeQFHN89f3LInC3cP4OulRYqm55ZER1kLMmDfI4jZMrZI0W8XuN2vCHqLWgy3VjxbS
NjbQrmILQ2JStefTprjeleA5vvbQv5gVYd6BoZ/d4SRtCzcSjvqE++8Y9tEbtO8zU6blLRqDnDJQ
QX1/y5lJTRVwSQ4azExDr7JBslBqdh0oe6qurPzvn0owBTK6zlsB457IOZH1NPGB4j60EUMCzgeE
e2L+0Pkk0M8TrN+Jyr3UJ07epyaPcdQFmAnDi7FNI9hFZhewBCNaSmyu9KdV/gHyAp77j0D1mEPf
TNJj86wZe0V41OH3Mwnez2kT/AXXTQMRF6Y+g04+QVCL8FFl/XGzLIG8yVPL6xp7eP6X63h7nmbi
+EBNkKNPP30gPOt9D2EhNLxo9TGMMgwokMK9jYyxy1Uiv1KJfeRyxPWhxAEFpUqHtvWNteemCF2P
G2v4pMKMqUQ/2aUP+ZrTt3oztM8NIrNhPPxqeghHedOJvNRImmXIrNlvqmJzJy90jkzjxuAUnbj9
5OFT1n6S31kQUbAyXZj6eLxHW2GI5nt1EPogQEfBSJCahUATmfxVeCi6rNfwaM9OJW8yu04T3bkV
9n2ejYI5b5wQqXK9fhlhlUGaffc8RI5KuftIzHja7onkS6REoVAb+IFW5Ip1QqvkdYUlga4oQXKG
vrgrMXGrGt9xP0m2phA4rQQNZgf/37NrA03olitnfxQKS/uRoSO5OIz3dMOu3BTef9hjk5cMjBBl
E7u5igarSlH7CBYyN3iXSiTkH7cVRJ9MYuPEdC/T88Ifhgiioh72D3Xy4ELiNUCgQG4kp9PWza4u
XGcTnOCNQ/sdUMp0SGuWUlRnwi4pVL0Uq1BFdy31JQCj6Hr0izBGXOEzUyHLS+15FMqkzFFBd9sY
0myxedBDOMI7qmS0Z6eD4MVcV8MrGT7EiXgJ4TeOo/pnKz1mImnvdXu4qF4Uq27SyqJ8aBni33Lh
EvJax+EXeXoJMZRVD9sRxcY3Fw78NHI2qS00gAa1CoU9F+q9nZc6Utu8gotDIQz0u42q1HG9/4Mc
diykdZIhJ1fHwQbI9QsB0+QnYDX1nIB/ZbIzKwP88kT8C2olOAHLhYe2gc48sQpd/uJ8Tg2cTtRk
WXNiVLqXjK9XegOuTrerc7gq4QVtiGRVxmM6KpR2og3KPmhoJV4QRSKn3Lw08HekPyz7FsM5wLvv
bAjcRdZMETTnlsptViLRYk23Ok6R4XcJQBRXNWZX8A60UQdzHpYAW8DR7fBr6gFbFPtYBgoDjv8p
IPMMdYZift0MquC/AblqrRfzgoR4YHHs3VpVU+jVoeUSPlikQA1TvnPkqLLBi/drWaalYd/HPx1y
FjSJkWv+kHfx+nAqoxYF+t1Jpceqt3NQa+EbX7Lq9jKal1LcOQmnZOWPtVAQKtF0wrCnEqDHUNRv
K1Sp8oKQAWpmtAEbv2W6i18Q4NZRx+MwQFgr3g7XnNIpFayVe7/S/rHM79N/g5RIApUxWRQaalfq
VZjM7L6kgx8FWYIaW9vNbmNWT5kIWPsZdEvp8nGPK2we85Wvf+kS18BQcWjog5hPDaCbMYNzkbsr
xNb0iC35XnddQGHHM7wKuaFaUYFjwm1PSz46YvdfAypBZJ/30FebwldKZJScuOj7Iw5mo7cMJnAh
I14PosHFpHPTjXDQrb0ZhjXuMpLA4F/7ymT6aJ1U2GFi9yJkv+kmDLaGiN0KFvJlfmOU6a/EAoJX
6NVMl0R3WuOFP0a1b5Q2utH/lL91i9Vsb1V2wapG0fZ0YRZsL14QrKKLmcMapbW0zdGINcdCt38Z
7q3QU8YIg4t3oaYOCBqK+mjhZanLLAFdLnfaCCq6WWfYVX8DcTPGa7HxX+qiuSnWyMIl9Ue0mNKG
dXOVIdG/OcljIhLXA264fGd7XIBJI4xdhtR6nuTqDgdt1kUR4FNAmy2Wh4U2wk98Ks2OTP6qFYSp
ukVVrWb04jSee1mFmWuKInS+JupHYUysNUK1X7FZxMQFrMPpJlA911iaYRUj18yCtZWXVwjxMUr2
Tiwqe0zcm3MYS5PAtyboI59RMLQGzi4uiHsTDe286f0Zw/7QXUB/RlrAUJ7T009XzXfLn412SnAp
Pa6gLr/vOFQBAw1t7hh13o6V7FHEsJWqWugpD9Z0hyAmQ4i8E28F9wYNYfmubEXXKZD/np0G+s1C
62rZ5Msn/xrpIBUUhL03lwEYyzxXFE92ftaPDA5n8h6iRRkVuPtOzyenQ9E3As+xjx/hLR2EkpaM
C7RruZmYXj5jTgrUJXWZJiApKdEXoj/0BpiGWk2Fd4RGOyt7P9If1Zm376J7A3U5rbn8Aj/5jinn
+D0XUvqcptJMuBJThDwqkVMg5/YrcqJgN/rkjTlOQjcZkTOzAengB7RuTHriREtJR+vw2gWjC0b0
xfFL7cOLy0uDGddpfVuFe2uJNvYFs96wqfiqlMn3YMfokLeiQOBMH6XsBq+hBItjnarzquyiHOGk
xap+5pfZaLCZzLfRMDnJzY8wQ8Ry3wgf9bENFmKk4Zt6VDT2FkFXeOE2CpCbCD8ughP+qcjumLpg
+71L9V2LnRL4a/bwHjVH0YWnNgm8mZnVinSPiYxqaO/emzLXM1Dy8t1xaPXfA81A1uY31uiJG6OX
APWr3nQf+t3HLcdMsUWDddD9Hvj01EmhiLCnyWEnyCq+QoZHbSDuwUevuOSGjGD9+xvMyIL/B3rT
E3zDhJjs1fz8oYsAZOkibGGP+5dfpJlWRF3zsE1cZzhf3BuQsLbkc/JJ54brYS4HmIulr/VSPNO7
DZhcygyK2J35IqaN2eTbR8+OEJn6FCbAZ9H68pDaOowGLSGqbtjheTnzIuSc8as/nmanCM1FZwXI
3Z9YZ+yObLg4Bif1C2ZM+ctSp5TocXJOyd5gwlFbGc6n3mmaoWszPzaR5RkdldzehagusVHXydag
KZefHwz5MxQID4/h28i3Y+VMF1jy131jnuqbQUG7Og+/ulUiLoEXKLNNgWit4cNtdgbTiK1NyHWV
OW/orhd4WwL23dte5QU7jfl+tFfe+z/9uBF+eiSfOnnHX15VYuoFfSLlo0ZNZEv5LqvwOInJTyNm
Kh9Fz0B9GQCCGwKMfyKA2i7GH8DM4ooT0i4O7gPEpsXyMroOctKeWwmHsmOjjWSWWaywR6w7zxEE
AowMJTPLVxHFsaxO7hlUnoNNeDKiVkEUMuLNFuqEYOGHU38N5xBowEpfNj0xi0F0t4siie0n28d4
GXn303gk8NxI9Kjk/gE4oFWBiNwk575X3OCXi3xP6tpz47F74NfLvtU2GyFAI/+59ngyXxPUg7DR
WFY9w5tqN9HLWkXXTSGUUW6qbVwYkBSy0QDbjI8B3TCNj45LYShBMM7zS3xxW26zKeYVo6mFklUV
snH/DE2AE1UY7Ifzo4Unl21MLZQKpZ8vExtzoGoUwBp2lbRrUgLIsNPYAwK9sUNrnEbTCr3P3bes
p1RxkhNImygguGdo/ZS5qTY+VFolQnNJzr/babfarQor6c4m7XnaC0beLQi81TSt5Ta/jcQlrV0b
7D99g0GyZR8H4SmzelXdZ9NolDLcz4oc5H2sOlk8XjH5adZtDDgsxSQDryh90Vw8RpYn7NGoOgdc
TCMcmUfxseCdotc635Ab7jDDThrMeNyvM2sbaT+Ft/oIsL9EvsIVXkcLRHuyuYg623hmV0RGWAE8
2ulFs+w2USBYNMV2PYfjKZEoQVAt0WvSv8HAF+wN9ILqX2Z1brMY2m7QUFMWHdqf9DkyOpdaAlM9
m6Qj7Aze3lWtb3jNZ9SkR3mQtcMNlImszlxBbh+ulwkgo3hw5wkCEV7ks5pGJcEd1EiX28bkTo/w
QIO43Dx6VJ4TNPLxF8xKlz1Zk/U5NLOHrdgWK6euyIpdbHurqdzgCX3ThBoscaz2i8fUoyBnCNEc
tenu1KRqECuq7xbSM3+kKsTnwoq9n6/x02GUSrRs7rVYqwAJKdhadIkhxyd8O/EbuHSA+4phvxBK
VtQx2zR/1BDhpfa4qqh6jWvBOtvlzLD+QNcg0f55nQxjbGMmp10zS9jDQDHXidiWsDvg7iOl9A7w
pRa1abelUUFM2G7Ebc2dU6TuGFmoRNTBUyUw/NSPWyUNxRuwqj/NN43uc/fuCy43PWWNfb60Z6VH
lxRc9G4421Z5s7bu0Zf6y7eyKyvwwkSZVOW8RB7V0HwGI49ZeqCYY70jiAADxeiXxCMkksFtNhsu
5Qpc3brD+Z75KI61/829sEkxQezGonCGvyez3RU3FNdUAhaPZWhgshVCwAF+/hHdfbSJ/V//qBHf
kHc4USfN4bj0HHSL3q0NMwgbdiCQpyvvRyukKs3d/br6q7XiNvHo5V1z6NeWbEsNHEi4x9UI5f3W
mZw2UKIn1IGheAZV2MK8pX8GJ5IFiJoVvF+XsrprKRY8gVi15hhNuZJafDR87T/3bkEnXfVaZAtV
BLK/iIqDZHR+UjKS6ynl6xuts1dgX9u92cSAC0MX54dIgRMTERFnLS/q1Wu1pjsUmOVasMYXOnZI
8dKpTFZAudrvf1axi+cFrrUSrVDsTuNMbLoTPuoi6pBD7W4TDAIDqj4yqmwfoIwhTr1tS2+N3pHP
VlxFVcDoVZYLMVgNAE4IaOmoyJ1xzwe46NeSBqBx7qvtYCHlPBGCrhU61+96gdowcyxE4EIzTIA+
zyfmKkhn8dV3tyAejuS5uQtlIwpaCzFFE6jKa2VNELpK2jZYgJyp7mb5kbeKc5ore5otTYH/QWN5
PBNybR1ELOeEQ08z1hJMK+jUIWcrSCvfbk2onFtlb4HSba5fRy9QSMrolQ5RNK4kZ+pnzq0ZzpsO
mFfRyLTUyBKb+X9XLn7U3A/KckdrZybnMdIWN9Gdtuar3fOrZu96Fo7QJk3vSoy0DBzUyeSkFSnh
cEDhpgI/j2C/Ojo7zhkN8n/N219vwqpFbD1XRw2Roi6jV8dsnTujhwzzp9nlCHW0CghFjKag/yqj
OsLUwRkllvO4peq5StnfMsQsgv6sxT+DsvCui+apOdUNtVvsDjUK4tm/010lwhwUnM9XRQBSz+hS
oatwdVl791nFZiR0ZIGD34KEoIzYDy6vj5aoC9RSc442aPNOtPeFcibxco81rqaytzeokqS7lPM7
BwOoXKPg1BSXrEMVD1gsg/h2GqsCg9elAeTNzBBJzASXRvjjcq1vGY6aNX6AuL92YZmD6Nva5ls3
fdgQxzuc1Yrg1gkSuCXZXEwm0gU6KVsDcT2Sd2CYvtv7LsFb1JaIUmOnmG+h2gnxVk4kfNa0WGf1
2KAcQfXmrCP38STrLo72ZWYuHAaKyW4e37x6CPGrPUyuyWUOc7+uWkfS7dcrtbyaHytft/zoUy5o
Q5ZCOg1iPCU8NZ0tfR9Jp5SjuYtsnCW9xBv9TU5hr9Y52cGBhyKnSoQ+nJLCu2b0qutYCak+REgZ
koGlg4yKlSmaqDYZO6/CTPm47u4yZ5Ebzr6xoshYn0nxniiDySJ0vjgNkZNrgzRz/RNI6AWeuYOy
9sgq+bikwiuXbVcZg2ghNE6aPJ5ZETECEas5YrzoA4bFU4fB3Q0BNTXR9cr14RKCPEIo1IqPWf/t
iGio9KbWen3uUwm4BxRk0/2NFV4Y5WNOGzhxzZKBv1+WiOu+8qh7uj6SBFo9b65lFrJP04nttfVk
OQunSw42WTJVXFt14ILnT7+xaqc4A6jaLIov9KbJpCl2XfzRR3UxVwxtKwAI9z9ZKDqWS8OzmuG9
bWvuN8Zv8pMgVeGoE72/cqQRtxIBT+ziYQi+byc7bRSWinX+eJ9C2sKMVAo5NuAUMrWqpXvN61jg
jyXr9fSqolwVa+cLJB6pn0LuqpeePLtPXeo4kQqVukMnUy80j+QBKiL6ODiVYLxQx0W6chvroQvi
HEQ+oMm2WL9u57E/RN3Dok4FCHiL2tXXtFV7ekzXEVubMUmStcmZDKvLJKXwZ+S+nb4MZ3KvaiLF
va4Tn/6dOzrm/UurJk47WKPBzMhccVL0cE2YDoyWCXT4ldvfHq8gFyBbj+cdc9lmNzItmCsxoez4
uXk/Vu5Mifs6S6u43mfFWhgo+RyEU4u0enVstqyhBLy2ZjPsEFLxZPlb80kJi10dZjQx/0h0qeMj
D7KMwHbCPKlY36e3n2vkshgDkugr18koRiPyKISrGBApV7WxzXSWyaAxYHDSV9QRJW/WSY1DBvWi
mlja5dsgs7lmQsLoHABS2MV5zYKo7aBXvdqN7707ThcvsZrumJyYFlgPC63NYMrtQs32WC8fl8+j
bghDKd/BWy++5VLrURnE7NbpU0FmULg+83gDLBgFzHip8DH06tYp8tRPQbCBF63JZp67mECj724n
lNFta7cBBoicijM4KSMbPpX3wMNGkgJ32XKGUxFdG/VfqXgJhAV+BvTJOJrPirwYomKb54CDTJcn
GYaat6jiobXbgcw6d8WtTFqM5Qc8RvBigiAMzvAbWCovGy3OdditK+4Yqd8FYHiQb5C7COu4pvtt
yadWQPyamQn5LFpq2CFe/5GBF+7pqOPc+BwDcJEIg0YO3Ca3O5r5JDelk0GqEmrMq6+JOJ/KgNc8
VOMTWVN0QOh71D1vqD5mxR6GwugFZ7Cfy68v08Gbochdx6iouSvnROuflt6G+VAe6hg+n5WpdLZF
UBPb91pEWeLoOVHzJSLflqm4aPkNvZuZHd3vrEkeEJ+AZRBKQd/qjY+5bqLSEjvpXvukHKjJP0+M
ATJvMbQ5dUBWAmr2M0CNqNFSdPDm8Wp0aSKf+aBzmVdDlaSeahewSU3aJC9RDFNM8PZwYYHZs1L9
ds6WDGzxjK6oF76S6Sk3itl9g6Lv4+8wV3UB6Vi11LA0VrgUW96cvTTO7itLln//knoozgClFm7w
yMC4D1lrNI79JK7rsPzECdIPniq6+/YZtRCUU/fAZ4Xgk2R5Us5Th4vMqjMjxx6m5Jy439oB19yo
65PO14syZyNGiMj2ZjG+NTVVM6bpVMjkZnhYQVs/ZRKr2k8t7TIV1MB0/BV3kdDhqloGK0Kr5ocH
+XCWBof+v+JtcHQGlvxRJ6siXhFKONB0ZOUXtO8r5qi0IsVMjfCust85Kqwbr1NnIRIc8sl8RojE
HLU8maZkqfGpAbuDV2VHAsrNtEX5Ob0qSYVeJLQNUL9Xi+Mts/XszL06uN0xZFFLjtqvk7f9zE5y
jABY94ZEVYRZZZZhkGVPHUdywCt3TSJ6wqeRnhnbqw0Csy8QXFOPMfWVf9bvJ6yjj/n93guDyMuh
I0VDWUQKUd4fHIPoBnEY6OUL8w/eWWCbG3i/4IUFd6lrn9wBjTRyp7FFzTTj5EoxZRSihJ/Cfq3E
RHiN4NPtqts9qbbw72qYfAm/pttgwFcH+9ijFtIK4LJquSFeKWT6/E+stzoRhMHKTzqpeub8W1T6
Q+njldNycxWhSOUFZpajgTwlOEF4I0JBd4TuQU2jCGX5yC8oeSCUR69me4LMo047XvKpOsGg0YUI
oXil/XkGeNW34XX4Y1cER4Vrt4gzRO3M15Q1iZ4OtgkX5+IUhw3oY4OIB1QnBsyTKCp86OWWMM5A
BRp6HiqoXPmb1Ile0aPHkpMGUr0N5zy/3e7SGRSZAdaqsu0DKuCt5jD6iMM3O/UwrKMEVA73w2jj
fReRJ/T+rcqsusbM4tYwR9uPMi3ZTsJ/kM0H2/MncXHChoBi1mkOTUfj6IVxKrLYHNRz+HlYDSOB
ZDZ6yDm7ZHtm3DxtTnkYXz5V236yaYw/crBNQqWuzAE5A4BWbZ0T6TBXDMUp8YxF1NNQbYSdm+Sq
vRBRIxGnTnMK8DQV0VHEKybrBSiqEnZrsHms7StQUuvTF9y10VuGRczVBQ3BSDdaSTQcEFL9nIXp
Z2F3v5856cepO8hc4LYdg1sR1RFxJ2yCoeu0MHmdCdr+uUdBYXjm+aG2k5Ba+b+kS4WRwONgqlJN
7LbJaB2V74t7C75iHYntl2BP5euEWjoITJEf2BMErCwDPl6/mW7THxHF/+jdSDgGmL7X6hHd5dwK
1FFH8uqBseRLNbQy5yIDyvK7XlNuEPD/RXQkqW0xt+Zrr4UyQ3wndrNgGO9fWnqNcsVaZlhEJWP7
7VDdkhTUZG7nCwiXezsMdEWB7CHMDTuZTun5HPu1s/M3r413wsGYSSZ1MENn7+MurQ+pAlK3Zn1p
BQBg3YwtVEJZW2/X0DtdEN45rdH8wCgUPXDBtrv+FRnRvCd2wJyqKRv03dd1ez+KmNDNChjFYHxh
q2hZcAz3BeJ15hNsMFKKLHbRTKzpOzdY5VY654SgjZwg4WWDqKcJb7GhH5aYBLLhJbfGTFUBx+rd
xs3S86m84830zvZMXQ6b5ym+M91eZ4t9Q1Usy9gKufs2cY7kTX7vamKGSya27syBvZFEFGkbhS23
S3Zv5sJIOrXhRnpS5lCGTUTsQcv1lPbqrczkdwMIRu78ZspGv5g/0Fdjt7NeUyUJvobCbOtIVh8G
wtifBz22snY5dN1nrpQ86JobfEcCjAAzoFOZj871h5GgV/p23jxMVwTAF1t7cmyJZaPx7eD2b6aR
U4d6tqeURb4G8Ce2+PqXP3NDlJOE/6FCEGsFxRf5C3CMD0KnySvrP6+tRsckbE5cev/fO9jdJ/7Z
85r9pdwDdHSMZr7nlbD8Bweg2Wgv3G1Tj1RIoIWcrOGbhMqO7B7UP6u+gGzu+LA0rzzn2IghiMmb
Q1dJpm7HLx75Wesbm8QtgqAY7c8MHjUCTBxmI131rV6D2tG2R8pNCNinLsEDRtsj6jZ/LJ822xKx
2yzAL8EzFbK0WWEUmzhcQ/FZDSPEmWsnWwvi/unj6badcqxn1fKXfnXP7AwnuQzlUHfFwKlzVb34
3qstMZY3E5ScPknq+kfWQP7HtdgjNup7u2kbchr6njgMbLFZEE6Qx2leoSM9DQsOQWLii5T0bnlw
Jwjn9QuQKptROjhEZok6+uNpnKwcAtqWKUBRS/K67e3hNtod/791EMN/ksA0XpcJ+9vdNM3NIPWm
IujbkDqS7VJQPiZooQYCCrrJErP7awTAuf30SKlsX/BItOp4HYWbEv920Byr/82IS4p/yFOHDfGB
ZWYxvW0I0estQstLrdiUt4Csewaq9BGHtnG3VYx4WPcHkMHLmEjKyER3yoKPZDqM9k2WwyvnrH63
tupLhGOPDV27plV/jhxUSBcgbN4a72Z+YhoTMDlZc91V3wMjthOJjiv7OrfrD78mOj9RNeqnGr4P
hSL7dxqP19ac63gmzI9KPRzlV7BXBMhaMtDaikdFTnyoMDDw/08Jjq4Z/yT4KtTDcbd8gyPiKtn6
IJgwoPIvVBxofLzlEyf1F7tBPqJpZr6Tg4cf4tyEh1YQlhPGUX7r3cX0eZFi90ooHGEjfmDOCdiH
ACb8KzexHcH+I8SKoNX4lmHMuN9B5UUwGe/OR4T+FjrdINx1yWMHA+l5SGvzyNk1/GxTKOG7DB/g
j5D85uc4oyZ24tJ8zdYkJE8PDb+TQiqzhndE/OWCRdGz6qRxjREa2PrSd+eE7U2CvkmD+YqTpmcb
74d2FQzbu4Rsxs6Flq3RnRIynr6Q0K3ySbZgKyAEpyeBvHBHLly2OOegsRH3D5y29QJ7YtCyWcc/
XLmmrC1K7LImC1Ho7a6MmcIL49ec0gnU7Y/4yxYkLe2NsAgApsStWCjHuYTbUVBC0m8n38s9qA4L
AztJeSPl2A0CME+NT6R+0cFU56zD+avSBy5rimOR83rPjJ7hchqP9S9LEDiTqO7LKWS1X6CSaPXt
x2ngEV5UE5m1R6gnvTsSYfm9T7nLUzhSsXbzUKqPgjIM/4SDQz53wZfMnCCkOMuTeVKA4DJKBy3a
4FvbKh+Zw3fG/TfCqmRzcTvOqKoxD4gFFHyCHQ+nj84+CrsNoXfN5hK2u/ZVrwFgQw/w4fbliCJV
ZnWdPq6dPU26s9f6w5SdXiHNChWzJYww7BLm+54Jd2HrBLp26L84PlTV4p8hthPTldyGfFpVwhxf
aixlVDqrp1jyXMu9asji+6wo1aHAfGUjCcGOt4TvwOpUK0uZKcD8TZJ+w90NMd8xGlX4aZtLFOkt
MAXYW+6N2JGNJ3PMW3dunGhWlLjtJDqRZUShiMTwtr4Rz8w7SHUZav/SN9oRd0qiCBd46vogfucb
UlxucDSGSjKHxbnIAvZtl458VMTtpr3P1eniNLFteAKlXLC6IYlHcMOVlMqYGMH9WkZF0V4r6mx5
ax0JPpfX+H8K3q8pgc+H2LNIJbp5OejEJ46eujYZ0jENvpW9qJYkWIMictN+QOJXx7NDDM6KBFrd
gXfCL3T2eD5yAu50C7AqUoNZux+hJgBjf3aplHzFcINKiItHhTc6LFCPBPfwRr4+e22RM8SHTq/7
3PN3hVB0pIV7onnXufRdH8HPcaEI2Yu0lLHCmku1BjkqFr3dIPhjgGSwKYqBpT7k0TlQz6uCmPyN
GBrHJhrreOHL/QYye5JRlzETc9QgkZ8pB68/o21XHfmim3yqGs0PRuQppDhuivQg+Wtb9fiY2Irv
Icxo2sP0O36/nShAz3kNhHEzhIEVcLXoWET75auUdmNMmpBTmURZLM4sgu72IcCf9LZOhRXtH24t
Gz7Hi+lZvVDPZXeM7NT9ADongTexBYuQuZMd502ORF/dRm3vOSN4A+zuvsWpznQGO68LDYi0UbxD
zDYVJqBJibDMqGbTH3EXCRDbyXFfYCLq9T7SDwQ3xPvzIfJjUeI7GDHzOYmVLYt3HnsVYuUnCWY9
JY86T9nVDMR06xngm3TlJ8m8tGv6w/AKws24PRi85Rj92bHLiKSZchq7jPqKn1bdIjKY8wefM1ol
MASHPKw23uv8rLz5MRrwe/EQWPXYGJYVHW0SEiILfaO4NaCZAfd7+eW0NqlcTM98ausShRR9wUtI
ZlFRtb9X60tMeT6oW9GZden8CoQ9zM9erWwgnxJHq4tVZ3PZgS0Dz91+tQ55kJebVaanEvLocJaT
5UH/rYx8MXzyNV3aIS5cmHbEgOd3IUt76l6RLDMLa9C3r6nrfisaGyST+OCyIGZme2HRzKC7fg8r
P+prc30AgscmYJdEjZQKmWVbRgAeN6ry8fLlKuKwNGarxvBahizHQqWQwhL2j8hADh+Z1kHvNrLA
cJF7aM44NHZ9k+mO/g9VF4jxE3a+scyh7GRDYq2gdeQFtuxYsDXKXm7Pxc1sGyVOqARVVPjn6ZmZ
6eHg1zZ1ESI3xertWgU1G+w8+IDZ1++dYSRU1xQMsTuDDAP8JwZ3bbffEkWvoO2oz2qblCKZl4Zn
lbjtPCjJi55JKNu+igeSBpvJIdcRjCPGg3NdfElNhI5E7shsquJitu27XN9OXjqyPqZFlapZQHZo
YgrRqPSJYvxsjYk0fjaxydAeodFzE6c5tnjAPXHtA7e+EShesvKlpatXFsuqf6sR5yL5FC4ZTEr0
5ERkx7hgF3pyv6O1JLeIwnmP8wL5rz8gmOE52Er9KgnEzoyeBKThs8+67nNesM1Uko/5DafaP9ug
ygCVEzHD+oTvhQtqCfyQWTBHQ4yv1B8YNpaUVuG+5QrcffYya0DxKkZmRFmNxsRODfG8ey4I5C8w
pmU9nZ4rAJ19fbQqf6p72F7X6zsupkkuzUenufPyrcb5YV/a9NRNjA0mz7b24PILShEKv4r5gDvs
ZJ5jfet/HPq1B8MfXRiInR8fSELVBZ8NJ1Rnm5fy/xN5VAQsWuD10YlmRsjhCcavmDyjT580+7S/
wCPKbKWAeTgZ3wm1KUiEGCRz7wdwFNojzjQY8taTSK7DvIAMyfLerVAL9Q+U7ku/v0z8G/LBG0CA
ISp7FRbCAURuhJUw8Phm7zs3i3iiGgJMPo1bS2niGsXYzdTbqNngoi00jX44saCWZwuclUFgbakk
QKpwvvCOGLTbCuylPmyrVBG8ZJ4VCYyf+oymk3v9Utvm23MlqyN+lCo8ls3Lbi3zfftQsk5CJ++r
Xks9MAZ+XGhXgwJOVvSg6+MdsooDP/+WNhGqGPd62sGYmOcAR+7Ay2BFvtu8uybAdJv/zxbFFuOr
/MA6HxAWpfKpewtegn44MMdlz91Cv8qRe0sMrvm26IabXMRqnFhhMB7+jBVoJrryF1anJLAzESTs
HXACCIDNqxJcILBZmiTq53/Y7WCTaIuRf+DJfYU1FlfQvn7sA70ErNpS14I6faG5uFqELr3RxvNy
m48YykRvfg2Ot7ROGrF1c/DgtSRTQTaMQe5HrEJurYvExf4m4ZV/nOplqm90FqqyrsaxUEHClaSh
M4tQ6wUyh9xMd6q0V7L+WRrKJ0nwhLMYW/L0B+pZpEvtqopG0/pYZmsxUZZxpn0a67H/W965Ib0e
ZG7IW16AkmMbYutfZTa/q2IFzhAKMIz58ZqgbFULtf1hTYk/2Ox/r1nxJL0qdDYWk6jnQ3MIL36m
xiwthYRC63opNmsG5lMZMrt5kp8rqqS978/eY9j7GT9FTjkFUkCfAT5ewFvEl3JFrroPc1j1Trvq
3beWdbFz+Cr3mqRUMHLOr0ZG2Mv9P1CMGRPWntPDh3L6My9PR1HzjG9dKqYN9Wvoo3Bl73PjqMRf
aa9vdk1AvDCQTCU2fSAcpv+wGGzlqBcCia+WRwR6P8+r/5CTTC+kvBlPFlqw7nFJrr9+5sJa5bsW
Kz5N1W+/80R1Wc+SJRX9Obz8jpVf92BqoHxEwJnRvikuIr5hOXifLncsNStpJUT+hT/Ie2kGbkys
Nfrv1l9Vwwxr8JCB876yWzfsIgHJtZjz2EF7uWpR37aEN2h54N+Nwi/h9aWqFq+W7Q6hLd5Sh4S6
wkNuOzoo25KJIWbFJtr4/P/S3eDo+Q54s5aVNCQXyFwT/R0VPxxM+eQx99+27QNq6rX7MU37xyuq
pn9udbBUP1NxzbHFQmoRZ49RYN7u54XxzmWgmpiediLHuSqrjBFXuHn9KYQ4zhTOttDU2hsPwH0O
7UdtCmFv57UxYj1ZJ7nRGJEwCgvZSexjDY0jFOkRC48EOpd24/h61iUjnEiSdtOfxYYLL7xGHKRt
68Rk6Ao9PzgaS2wh35v6KSrw+SA14h+HJtROlzIhEO8Qt8y7fOUxGZ1e+Hy5HP9otCkOc4zsL0Ce
bcnbIML4aDfA1T8ldWJnnPvEss3p3GZsMURUhhhqoK+7R4+lcDQeOAckPr9cTQQIlFrs/C7kEU5G
AluiMtrgp2t/HQqkiLRuvjaZzLlWvvgfYOEybJx3HbzeqSOgmX/Hr6/qpvMxsl+IxAjOq8bSSJPd
dCmK0N0jPcpsvYTuDwXEGapwD4TrzwwgaFdqTe9l5rd2nk545sNFH59WvnxMW4g5HFFGKtT/EetX
fx5hI8nfphUAo4DPhpu51AgOHLiwVBj46jQXi2Cl8yfjZrwRk4n4aTuJ0tQUyBfL5iundu44r6or
md7GCrgx3M0OQLrD/V3DRQIbYQ/gLQ/ntvQjiSWvpde26xhnOj49I2pHF8HOkKi9geU/2pJCsq16
4ttLEj1j+1dwtIq1UzbMvsKPwT0o+BZFZSfzkrpf/t5i3oTFkPgtBN25rmbE4IQVYRQbhxggbyMv
MjsJrRID7zfKApO5TofvFAnd86H16Xb8F22SHrxQ92R8ZJj8qdBF8haHCzY1Wef21B8GbQBrBu7h
wEyCmFEy/pohLeZsA5BYY++psr2Xv5SRWPjHIliqihxAvxKzUL27qACFORCBJ10hq/n3rG0WKcOv
/S/pj5kZBJJrjBM1h5LmxhiXyVZFcNk8gIgAnz2bqhlEh8k9gXDzpPnHP7hh92kEQpIr5HVhDSUH
dG/TmZ+GHbN2OFZp3YdIwgU2Orq0RCMsaJbSRXgf2lrO1eGlpOZrsoQ2i70BCrOfn1fNhoK7X+C6
hxnaU5WJb7p1MiTx3fYTY+TrGNWD6uvL1Q+RGaeGzwYsRhOWx7kmyKcyJ1/iVRxHgsCOo0ciIz99
geWnZCsXevLDMQ50GeNpvvTgJScqUegf9LopO62lz12m6/6aDdXpuyuKkkII01Q/3F44iLzRCbXa
suTnr1HAjcZ2+KIK0tmqVTydSdjbx98/FM6skQsbCyXg5UBSEvHhtoSUt2UMSmisz3lYNG8W+5vY
cDjRWATuUNXwoidDlo6uqfKh6T8tCJ2VUXE+gbPhM6G9DzW3FR0z4lPJdP8iD9JvPbrfbUohFFyd
SH3ZhpSzH0UKZrR40wUzgFg+EyBcShlFUbC9yPInFCDAN7ZkN7VSUNRWcyE6Thar9lL0PzzVM8uH
bUVP6MbENOqSE0OJwWwxKdluJuWiTRarQ8qsco3KDcfKG70mBbNuXnhEDrdBtmS+jww45Gjaayhx
5mY00x1o35Dpl1evyJXBqU6WaLnfMqCkzmJF90mDlE5J7T1wDRVCPkpkbyeOTEelx+UG/qOsiy3d
lHjlCD2tjGrNvdQHTCixZlde+OFpLWgZrN5RX9cYurq9x7bC90hpN5a6Y43mBVM9Gtdwo3gyzO5G
P4YKnn3veQY5UIWd9BXE2f7WOV8UUTlR9024B/M/XbqXMDfzwPxzxJGUftS9wcNDifYGJ+N6dLy5
ydAR77085h9Y+iOwQhOQ7c/hu6bvfFNSVZDS+ZryX+hipcbmED6phH0u0b3wVOCRnmUQ6OyMmGEg
vputvPkpPbuwX2E5GAge4dK/6Blc5b2iKMI0rB1QFjtLUXUzHjvtTwqYK9PjnizOTfdivCGoV6bt
DExmeVtEmdoQLJub20nbplTwIN8TNONGEXnhHXO96b+KLTlkOfrOBJUGKwx4CgDgNSEjEwSHTJrJ
/3r9CHFKzrdrE07Rm6yAVRA9ak1kmYXhu6uq5RfLHQZu7f+rweG6q0SfcrHz1wqek9Tju0Om+lgT
qSC6U1OL8NjTKIRkZ1HMt9FmyAqHDXpA/3nTVUuJTnEZLxYIOGrjb809Gr1iBJ08uu45VHLUemen
ky6PygCdBKcwvhR9M2bD0+rydG9eriq1NTT3JbLzDSMu7xW6uAQbrpIlboaL68c5MiemB4C2JPVK
5nklATrstZApzoqh91feIYj9nAZEf3PvrknUKt9Yf/H1bK7A6ZR/jQQp57UIuZQU9Dx630g+dcs/
OOVskFUye8nE945nk5HjzHO6vkl9wXLJPDYvboegtnuXXvbLSo8yHaHN4r0tBZRvYQFT6McKSbon
60wCNo7iEbslJsxhXPuEhPnLpgLg+6HU5Q2qgj80pou3oVhopZR/Qs0gy5TtJMpgbP1Qh5Z23cgA
VDaDo9NxLrOg84pLzoHUGLCzCCFjto49l6ApeWgRrL6sdLtu71EUKRKt/FqTk/HHxK/7FDLABcJv
w5xgpgUn076YLkRBWsyxdE7qdFhSEQfPwKPT3MGEPzJDuTyRjEEdF37JrTriVxhPzZ5qFBfms3PP
6lUCqf6W0EzFYoDTRZiV0WEGVvbDbH7UQhlYwhI5FFswLzF89VlySf4O1ndRNeKQKFCqhbeIPEgQ
T148xRApIZ78dY2AmlVmAwqib7V+1KTOExd8EvYt5qPK0oklKDZ6OLVziFE/AJlHh5aqegUn3s5u
xTcqKNCK73/aya4DCmAGG8Lrw9anXucTwB/htISUtiQvPY3k7RqYm8yMvCn5fSS04ryf1b78F61x
Oqa+qveNmz+5reWzMNQPHprI1FkP8OMUJNX0+3rGl5qEK9tefRBfSrLWWafkikzRETu0rgs7ljn2
o+l/DrtXEyeTqkoyozcWsc2l5lCL5DrYNSh+yNeqHsNJqOu6EAEA5q5vooGayH+jj0BOyw5jz0sY
fX5RBFB1ZsqC28Bxb+us6HitgDHkAmrEmsgPV2ypFS2rLNPhN2S8hftvc6YDb8plbmTEBrCR7C+7
87C66F0tv4XYSoOYZQZunOt8llNIvs5/sOKet0myETUvi0J4byRi4GhF6lo9qQ3jnLAlJOuWAOVY
OMg1sfdoLv57NFNTPVp6dBnERVhiPmJnZlsBcixnncEsq56HqeE5UjfXaTB+Kqjo+gxglWhp5Gqh
bp2DkZVDfpqn5/yV1XUGy+sS66foCu5nAiPdvlEztMMR3nBun5f1+y/dUVTGMBHKDeIp/0NsA+we
C3Yzmf73jpsl4r0oWK04p9SZJPb+osWnRUT7e9c7inch+wz9yK+7wnKiA+VqF1jRRp6sSqB48dnP
zojRNbPPoqd+k+GxG2HxixeRF+HPLpWmHxdaduE4I8uWkWML+Vu229/IysyUJQ/RX3mrQy9HiEVY
mLdcoz7xcSFBtKB6WRmFai+WoTyMVeepDnhTZbpPHtkgmBt5lFxl1zv6KjNFWs7ahiUzpYQF7Moi
Fw0QlfUq+2p+pKiBuEtK3DOYqTMYPRMGXG7HrU/robaffJAQNCWUL/Z+pzDtjXk2nT+9qyf36V9e
qRduEjOG/zw7PNSlZ5575yvbIZLnQ85yecMQVJw4rjn7SaT+t9XJAITTe5GuNO9iwTGkQBRUcZOC
NXdzFexhdYyAUAf/69KeIr0h/DtZ8Uchlk+XU35dzcG8dSZ5XFaQ3GPCUk+uUV0MBuWtzqqPQzrq
S8KpC/CVXnHzaS7MukWd/Gp0/cEkBuGFCPmXiHIpeNFC+UO8lJeP3JfszB0rwI3/X82hBUdzCaWj
2/93FeSi4Lr24+gj+Mx+vyjkGLVZctc6HUuY1FDW8htc8Wed2PkXPELpURAEE9lt7JYxK6XByoZL
Tz8zg/+72hOXDOdSJ5JcOravyWeLeutCD7D4deV4Wgjn6l9SvWr2ueO1YV+s7t/hMDqr06cDC+MT
GDSsWSnDrqMDmYS5NteqwvMG199GvTfXXDKi2bWE8FgG+EDgX2xYj4xC5Gsbt/tOvuZ7BSJv+yzm
NEb8TrV9TGMCrRatjRNshFL0loOOUj32eXur/61FVTsPOAPLGTomWkBx22Z94XDjeW4UBJAsVT+M
CnexRyVrJZ71m1F3OmwyjluOJBeTDODGLA22b7eE8dg30sCekq27DVDGwCLaWqmdhtNw821mJmDF
zySK4S/3qJ7fKO/01Jz0j/yjR3XrTnxr8df2HWrh4hIFutT+CLVSyYHWUx80NmrHlU+eFTc/LUvA
bdPkCPsTnE6coiSutdIkBO0bOISfxoplBbPV2xjPrAwDqAhuyOhrgJ6fTyEMzD++yvEr8cN66NNH
pNRBhd/sZDtCWwz/QYBWsJsKtpNmxcoVLjGmUa9anDRH514UxZv51fD1feD4dWrntaIfxagLxU8U
gYT/yKDhNwJgzC5S5bJ/4iTbzt0+ZDWXEUM3rC6+JotcdlGSyoa87MdAeDSPh9xl7B3XCjfp68Lq
msTnnyhthZd8oKStnXW2psl7sCAXtdGYKp7I1x5Vt0OncmspXeEGDkRmBX1XLDpVZqjUW52j1m3C
xF/HrxiwrfRruAZb7k9bla0ryHjgNwEpbiiI/LotRyqhF+Z/p44KVv9rg4k2CW815U5i7e0Na8Pc
CkY9nzBFycghzXMO8/v/xAGAkHh97NYvpeqWSpo56ByWC4Uqten9wNQ8tuFpKjggjix2JdwFjx9O
8VzktEulxT01PZ0bU+LonAwP7OY/Y+5MgtUaobMt2MuCVZqXaOk/D2/1gwsHXNJXufLTRUxt5GOY
/DlWD0MCR/gHYQfgR9NR8vMVQicy/OVmOwuRlxwh/1ihe1SMIop4TQKCy1vtlqi9+1r4ZWO7DgXC
wHar0uUQQjuiel+hQyXf84d7SFdXddXGuBjolDJf9kQ7VgM4kV/v7o6aB2wJyWWt3gNclorFgwWf
Eyszd/ukDJtmzOatKMTb++EDmRv3bPH76pGBE1kDDSBcn1XF4c1CrTqI/xiXqQ3RHz+Jr2R5CHyQ
QhCe3Ztbn6k39Wk1utaXgPBDmk/VZiv1ZtDI9Lt1xBGmMMh9DirIHFCmhHj4ua1xpvEn7CCFaoia
4QlA3jtEToUN2r6h/43vpYID9dCEGB7BU+7cbTWlfmbWH4ZHbzvl/k0HUwIePTwwZDqGIsmZTIOi
ALniRk4QY2JGczp15igXRVTBbO7bU9ZY2rmQgsB3qx0spHgNiL7hTjOYK8N1o/gPWgu8S5LZiVfF
WQ27McCq2FRYHJ3gs5UeAws9MOZpG0W70bZW/u4882HzGkbpIxDdP1CRuJSImNzWlAKnca8sZVY8
h0lGRswkYjDZBnreQx4W9A+n0ZopmYQe8w3+U0HbKfu4b+1+7hR52Ake96dv3Ui0wvYwDFjrF+Yy
vsSuZ6Ns/E1jnPTL2Z4ygHf/0pwZXQ+SA2WcWgPzNtaSJ64TbtV8+lCMMnadVFiQrtEpdS+ks2kQ
FYzULecv76CNtTrLG+zuCElhaR2slQVensxxk4TJKlkLXcVy0A0+dvEsdgxuA9dHiIbQ5l1LGXmm
3iN7JfwjTPwVFtFSkZdznHPx/0h3v6CnwWiBQb1XQyjsdDRMetEYZJHNQxGpIZvbU1dNR1/G+zpk
98u0mUNuhMQs6iJUGBQ8dI5BGryYcAHCyjRS9Me5Czq2Va3eZpsDK35SI4G6L7mkg5JaB4L+a5L3
TC5YTZL1UUaVB3g09Ns7rDj5tXX1cJFt8fewvl5zGw9LKoQWjTi4QXQoBWhte/FOBjPvlEi4sIb+
DaQKwvvoJiAwP01UUrsJpCQ2m9vl8f9qiQ9NaxjfTKsGyLGGOjM2kT0YGDJ9sYdwohxOGAthr2/w
JGYn5DNcG72EOjBy7Y3qBMuYmoTfnyAXdttD///Ks8uU5ODUXJzXqZ118vgFyCkwKQsiMfcRURPe
juuYb/13N+yvxQyao+tmANTfKEr69os+TMyB9Sq3KydPPZXcdS5uRfnI1zUlwK563C51VwUQ8CVS
z97tZvPZC96+xtxDsZ99kNGtSI0rHuBGBzS+Wbwzjk0L9aieeBmkSdrd1X/+2NmYxr5a+9XQaxbI
p6M/DR3f6sCQou67/8dgOaQpS5JrQpJTcByIKOZUqilySTgjRk7bJpYCRebmOTCe2/chNjaTm+zG
YndlPUsheE/3BFfGNtjsgyTsb2ngZujI2M8A25U/NL6Zzrlh5S0qdDb9CKxRq2I6fXNJmq56Z31+
0vhyBWlyo8A6+X6jkulaQnFAi23ccDOhUav9olSO3APmADz3VO3gEZ6pm3iShg9SJsgirt1MLU7U
YjcUdj1EdTXakLWoYazPDPud5BJ1vgsZuwXqB9XDNuVCQVX5YjPXDkjYKBo0z5NRW7nqTkpFZEeh
rEb602NLMMSbn1PGXDQe9UONayT5fa680WOywSPoYQzV4pycyqCym8BnLhuFTvg0Ttz+hYzdlGkq
ezdZEZi9EX9j+q2w69X8oR6eXhKQgG0elkQU7lhQeWUlCqLYea66ppH7nh1uZ9arCPUoNbTfHW8x
m1rGGRs086jdFLfOlUaIKIeJo2/8LNXV0zdDXBmzOmDQW+CY/NvrK9EPRj8t7Ecq5ZogXRFNmo21
YW3hCe4AQzatHd9dFgm1fhUKf0J+zqIQbq2BKUsa5CYgEG5JkqjEkdCvHZfsoXqk+JiDVALKqjCs
AZzI3vl/4EwHmtPqNLRjfSSpf0umcqR/1XZ5tYUoPb6i8hrLaoXYH4XGYH8LBDSterjsbx9I5d7q
5JqijzKT/ClT97yKSePdfvMqAanVyoPaoP8iOXIwrY/3qhmd7Tfuu3VBAY+qIdPQidP1gnU7egLC
T7CSzM6DEr1hK1D7UZX/sJ+x3mVKBcQQpcWMSMg/68Vg2Kwa5Y88LfEdvFhmsijKMMXDPpx6qi1H
uG7YcDrzMtPO0ibOtGg+uyR5yBncsWUVD86CpKBKle8nVFGxRt7e7xLhY+cqJfwRg9xZcfYZ/Lqp
xAr7PUIDBoD7pEZKMMxIKexSEmtfR5pZ29DOmtNdTV0Emsiqf4mwskKGSfuvSl5ezj63+ZQ5bcij
dKofrSFQT0iKUcbwQh2erIARPfwauEeLIRt2cWPCfFhu87/4zmvQFDlrAT9IeYg0UhC01DKu8fPC
bhH5qiXt2CIx32eTmnPGSyZyHp83LK3y+TtddGVwXtwRBW840EmO2QEYKPTFw6Xy/LXj6WFsOUxy
Pu3De5LApSpk4OQOrmhWF2vIzFwUDROwvjACL+GFyTr6E3ZYGF/oVc7fQhfBVjsnP9deT85M0KBx
R8X1VMP83hEKhOolbuVf1WBSG15JOj/HmMkHTcom1o8iSIrB09F/2gR9E3uemo543/7sIzyazivR
KKOfrkaGvGjUZ5AUS1mza+rMBbmcJbAgl1LXU5cwG5jOpGU/Yi0kR5DIdOi37EATnQTih2xZpbOk
3jdY6XEuuhEWLftG7xEftM+SGCYqxK41OwNyyfzpSymvxcgli10bGuRNDce8STaRmhykseWi2mZm
e4dz1vbsWU5PaNO/gICPN0qBg2jWZYvra0hdOJU1OEvSPRy6vszXcUH2QALJdwEt5qHWC8r/LhHb
gWQn133WM1PuFjV/UYf92bm6sbLSv2U7v367hk0P9foeuC8iEzPD+S+vwC2wCFktKMPlkGrwXtjV
5QMiNnElf3tE9u1pd+Ijs65ttE9kT4FAHDr0VlIxtm8DcCMk5OqrHTu1sFrsiRV+Oxe0p1kHbFxr
XjZTBbgzMAD/+zwqYU6AN19qJAxx8sDJfgTwLMIrXrDyJxalgE54QrvP+Vopvja088oMvHeZ1jcj
kqaw9DUVCGUUQHCUgKTy8ke5WsHnItwf0cEdQj15zToZ7C/s/pqA3XzDwQAwJOOPRCW3h2o94llf
IfmXEl1uO8RCeOHNPZu5ob0aZ3IYRXwq6fpLbIpsMJEbMHEfWIMdh2x4f3q73Siyep4feiB6Dzc9
N3IvtHTj4eDIhRm4L8aoNfNtnH60Wu7c5HE3PTbXLB6qI7QfvOtaQfAcHEfVDghoRG1kDzmyjYFj
e5AeMwks1RmEmPvVZ4u28IoY32DJXrcnQA0iWQ74R4ZsKjmqlyEw5UcbNhW5ZO9vHPzvbJcdqsxo
hGJnyux7ij/4vX+v0o0eV6cFWxgIaNSxxwGAOksjUmr+3u2SjDk9r3D4K8X0Xu88YBxeIZDPhZ5A
DgfPMSPGCJFVcvFgCKjypqURF7aiHcJXzceQMmGJf/l0CZpA6bMjQun7S0rU8e4xpNRX6M2En1TX
JT1A9cqe1ApU+IkYN7V+KeRpChWBRnO/UXMkx8cOB00XRhQLXfV4OqD705TaU1BZw9iYL47mIIwY
Ye6XhOUG+XGZQfONu5Rr9EtWTzVLrKPRRom45DKViYEPX4R89IALQ7wmUueFpMQlIiV/2x6P/Lls
0IyrNNDdNLElM9cI9ka2pox15doxFYqSa7tctNc7aLGc0cbhlEqE7BNPRMVWLQAHxsp1RiNIsCY8
wHLil6YCG8z6wSqtPxI1tgTFech01isnEWaYskAHEmYUpaT+4ofHrGIFZA74Cy56TA65pQvv0qhg
+imgy/aX3uJiSGx2IYKq0t9pETJ5WiBZF9sFRL2rPGdy57ge7o1FGlKTW+7nNlSvg+aSgcG3q2EC
ojRFk9q39nM/FPpDoW17XFtEcjUy3iTp54hJ5K2oORmoRrIzt8nUmXrLH2OvA26weT8DiivdI5ya
2I1F5hpLVdsbQwq6i9z49WvDd9OBWjCPearoKHo7Q9MWQL59GyttJsH4Ew5YOUDW1bsqTpQcC1tx
9vkWS56GdFzDweOFjhc3ORqJ68/wFgjOMTANfq0FYheV6NilZKUZwdElDf+Y2TsNnK6TJzkYOeC4
QxkhG95SC7yPzDd9cAFuDvdXZi2QJlBm1DdcSpoIbuw/Q62rgtoaOvxH0hWnQY1IX/zvAjsDzwRR
VtyL+O/pK8QjjBPm24iVRuhFDeen33ohofB0hjI6FDq+AaAFqOWxC9pm3o16OryVVSUVsyiQ5EtA
J/9JjL/z3ZMtfc4EMeR0QT0zFPe8Ly5TSVgP5qUHXdQqjusBFfYa9n5OJMxWD/8/jPcwQIA8D4Go
zVsnakwDCSC2ng8Je+BM6wcv24K3UU8yBnA3h6qRnPWSKDE3kWT60ehb7QC58ZGbt1dXxSf1t2jK
qkE8d0Dv7tyhn1TlKVwmz/aCqLPXpnui35Hte0YEIq1rYonMbdDylkgddHAicDn6jppWo8fGbQXu
fBbSZbu3LdVZ2Ta3MJac2/hQWwglcRL/UPELCWEBApnLsyPCx/Hd0EpwSA5u7vc+DkqAi14Kjqzc
h+hPmKIseDy9udZoj3hgbqjZKZ6lI0E9J+YHsFc0TZcsn/S41MSLzRDW1LhVhKzx6N2nr6e1oA8j
2cgr7GMpYx4q3WFKVA1rvx9dpAwLyVv6WSvW1XMDRFjc5HKb0kgyN4ciNOs7X7/TTRd0lCvr0lV8
DOrzs12m8GsuQcdZHpjILHIU+nvCcnPTzaFu9Ptnjy5bIche/nAuVEcYDvL9/AbTHT0egC/uvktC
0MVFj3knWS3keMFvricwcN1mU1xi3G+RcNavKyGtv0DPUqAk9/p/petrMXvnhlZ9iZeQSUPnJgg2
4nZFMkXp19BTgCHSjDZai03tzMPwgW97Z42+crTqRmeoUbBwn/QzOlr8ehY7crRxslRvWrrptvZV
XYRK3xWRrT5uuXRJMHGf0p2UPfuvvVOt3glvYIPeO9z9IYSEa5L7XhUoMvbcJG12eMZ/vhrGJUE/
qZYhAYp/yfDQWPMW5W31gGV+v4jbvCcQ+aNTXKwqIb1krDS910Q68prRXLjHuc17DoIIfoxtyWjC
E3LOplLJf1Zrakq8A50fVbKcR64rH+FYE/5x2GucRbRpP0MXSFoPlziWY0iyjT9I16dOj9atVjWh
Y99qHv/YM2jxWhOnCh5XjhMgxZEWB3OawjmSxjDSFvBzlIhIuazUfhvg/OP/m1AIQ6VyHJlMNcF2
p8pexwGQHJHvuNI1PSsPx0wtYEvW9Cur+yt4PziEkjr2w0SF6TyHvOoV6/k1un4CT7TGtSuT+HeW
6CDmlj8qTgjLXXHiqgunHLXJ5XA+gkk1MHp2tuSgjdYuNALhQ53UAr/0jjQVqcQBwHj4ILLWR5Bo
NSKF0ns9gKhMx9RHwQJwiDk9k8YaLfBuySPVrcIy6KLvw6ekuDvU6K62jpbtUcbj0u/qNx27L1kF
MI8KjkVS4QFdKXxzr6kWW+YTI9GlZX87H088nyRK/S9tC5Qnw4tTu8wPMHCo3QFknZ5Aec39dCLw
4AAnGyhhqSZFq6mNkgwSy0b3U+DT/c9FjmJfxYQaPTcq0l9eHv4slSY9ES2mYbrviZLdKjNGeDNZ
5ahq85j18KRn16tPPvjIGFfOJOUqw6MD81SxYsS6nEvSM9BSrj5uVfiFBX1vCNRgUZZpGAruSBK0
7feIppOrcuqmJ1Xk7xL7KU9I9sargtsVvhBCfJWr77dL7DANf5HE94Rz200uYemMt93dcaYRzsS7
KRxnwrWdJh73cmrTKneQP5S5lqgvq6SotFyrFxbObgq9wUHUwGIjsPMOBTBG/j1+xXPLKr/KWfeS
qCWQRD2szq5R/xzBDMPaJYiFHtL8tir/Qnl67S3rugWgd6HymaaZm42yHom9JlgSUeYbuWEjJ2ji
CEdAK0gVOghlBU6zJ41zgCPrYMAyqjjWXFGzB3FQvpuIWqU+GsxCR9HwvO0j+P8000Fz56G0LQW8
JUBQ/rhByopxMGYu9jP3I20QjQDbw6grktsXv5nSIWjDmPaMbWnr+fEUzcI5GCH0bi4JVATuyrTb
lYowPtROadcjsxk0t1w0J8we+DIwZ4MN+XJ+RyqQ229CVlBtxzyDdTEBJDg+Jzref7YjKnSf+tse
7fdt3ZxxXYb4SA9fYX7FnS9EDMyWB0agj33hs2YOg9Lt65UPixQdJjd/hb9xA1sfJZsCeAdN+Gl5
SoB0WOt8lcjKTI/j3kyWp/b92iHCjnr34Mmsbu5N/7TtiDGU1Fw3nwqwxLWpiGe5lT0pP7rMlRah
K5gGWkHrDyIU9T30CFWuqBZ663c3EI5nADzQBvEOhAhNx2G+gf2Q5gaI8qvrBHi7HOcfMKa0sbGo
iL8KucRMpXpbmrii6CaOaU1gpgAKSpEHEpRwud1VBBCUC2DtPyxTDNa3seaIrjAQahpTBSirelH4
ryACo8xVqBcsuA4S+w9i2807THdzhAxsla1GfaNQ8Zw+vkAaNWAeqmtF2XFK2Cp/Zvjm1mfITapL
04zpSJwzuOcVzll1B5oWIiKSPYCeWlN0AFHXFbcNK/SF33HwnrBAFwwg8642S3FR9i0ifQU4oEO5
y7YL7tWCPdUjIhGHwvbjNdoDs7yz0N+aVkY6vAvJQE7cUyiHaQiAftemN7V2PPVKUVSOrboVm7gS
mrqcb/eYB/d4fUbz6hI5Ny5ui18oJfwLaoGySh1RfcrECellTdSIxoIJRSZX68T55K0xKS4zlqvI
V3XCbTX1tpntMnrn1kE04ReoYZVhhZr9GHNqTh1xO4CKARs/1mmKG9SgDtDOsYU5feYLCLbsgmsu
yd0eE2DxozdsCF109PAGdDN5v+4MPr04X/XwhkMrFowJAnSbmgt86mFxrX/Kz8YbpNrPgvU9/vYn
5fs4UpBWzWAKyptJiVut6dspdwX12pvyvwbDxFOGl2fQIu9cNB6SZLvKnATDZjv1Ts5Zy5dHpJYR
NvM8LNQa/W3tCIJb6k98nLEVRi7h4hxNJHAHeeu7J9pCrwHExrmklM7HKYrJJ0kmSv2dsgdO3ehU
jFwFpcH/A5BKGG9vVI3g9/Yl52Bed1dwe5Kup+vg23VjPH90WOng5rZN+a+bGDGD90jAtFLfKd0Y
RAOGm40ATwbiHYs5E1CU6mP80fQNZHZP2xwCnEo+Ce8lM3OHipAURjCMFhhDUEZC1umz8fuEWBI4
WDQxL0dHnnbO8reveTVRj6PUZ0wC1ElCIRzsaw2s1vSclh0iaNNo4X2UCFbNaemf+3vi1M9+Z5BO
zw5CBgfiHjl6e/aKknnQ2L6eAZ3GhUi8w6pAdbhG6vExk6ZjoTPE/n9Rcr9zuv6rKbS7Oi5Sibv0
KduXDiFhycDzzP4KOrN51xbkDe9B06m1/KvNsuLbYN+Z3bKsgxj8SvkDudRXaKKQYvtv2gtjdBNZ
lVypaNlXDR98hiUpA24Lc1LxX3+vrZwisAzo0Zf5UKs5kxnFXIi74mL0rNh6NUc3kJnftwYLnJuE
747xQxtv4KHfKdWqlOaENRHQhCFQTHzp7l+3IfdGItikBy2rQ0+iQmk8aa2XjfZL2hZEWcReF0Wd
RiALNfgmeIM4xTcVYt+pBMDrncpZVPG0bZZb1NqZi47TuGJhkkA3wKahsYGTXu+PLYrsNwtFwFLK
Hg/9SOSVEw2Tf5dSNAjHTdRxMmmvJXTFCjsiRK9g/j9xMTsYEeSRwjkIP18mOeGzDh1yDhbEl8Dp
NF1mdFoUvm0AWz7jF+boDmeoeCjELG4OiJ7gDZYz10kym33CyTKY/F2LMhwVAfZJkCuw3WtAM/UJ
a93ZzQuiT6j+/DA4ouwk7VMVWogLxw7jIMvXpBf/mUT3G7tUYRIAbAYZlVYT6UzBUBU4nC3PUYaD
I0asuyrpOodGtbkStyKbCjo7MLW+x9iCWZIk/lWSLSqGfo2QfsK2gySqBNIkC/KzK1p7X+AVW48+
i7d+IppFxcQUC/AeX08N4H227w4ZKgWIK2kP2B+4u9yN9OaKnP0c673oS0kljOvZuWBmTM7+G+jQ
LFAMShFsQIr5VDLAnFV9N2if/8FDp7y2dQ9CvuKS2IiSD9ZG9mHHfhOzjYE94JUWroMPi6sC7gSe
p/FJ03ELeYF/HhHwNRD7B8o+3mNeuD2xeLTPBqloUZrGZ/JibVIfsci+neJOULAcEuVGHnd3qP26
std/v+keJDNrgM9vJjaZu4ydPAon/PGtuLwB8q3DYmnYiR8Xk44fH7DbCfCySLjNDHzlJzVSvfeh
iafjwLOANANNx3sMCO5J+BfSBliaMt87I6SnSg17O0NxmEAS/SQUZ4vmsSjIHg5HYkdpauTFKAd1
cn8j9kDuM46ZVIiaAU8uX8zQ/N8YmfNb0zdYdEtaIOTlkcjBw2/0X8ScJmxgsxVEWHO4HQ7Z6Ezn
v0y6KR5VY0c689NNpLcbWLkk0LcL1etaW/edrziJMEDxRdkNCuEYkjRlKfLyL/5o3v+BT1NgNCOs
VOJsy2H4pqL5yfmVWikYH/1GwmAKU6OYCuxtJfLcD8YEbGbrqaYk5mY9AeACxHepCuQsCXb3MLcR
7tFDmAWdDQ4bluu7HVoJVa2jXqrTVhbbAZR7lCr+9HrHabbnjICgC8w3vbzNjdqI9GkryjIFORIP
TM2r3zCcUtKyUrxNeZkr4CDIzam+SiENoo0RzVbYoUMOgXMv//mxvUUvNm0u1gGBbO6IfYeEyHL5
g9TZCVmPia6Dt330WBSLmPdNOmeg9FvNo6Q1NWgAFR893WHf1b99Wn414HfdhLHJWnlxgL0d2wzm
q9hzoyFnBEeT1r2jM3bu/++0RhQlutCPnxzi1uTQgX52Ylln4F4LHJArp4MX5D1FD8yq5SjFG861
OEaWdc6XdatqGXts3vNnyJ556ph8n12KnhAhS3/6Dr9Q0IFUXaG/miir1C5amEJKZtO329+wxlQQ
FzkXsUDPnk4gOjoIWz5NI4R2fq19OfylLY6H8p4rx1CfoYM647D0ToQiESCJEoawzlY3Ff4/gNir
2AKhMvYQ1WdEoGzbGrSfkiZ8xsPcQ5FPjS3KVmnDOqyRZXU8DnbIYPzkIusZttvx/lPYT1EcQ2Z6
5gah3wn66RBZKUqUJ1Ix5lTbi1oTemFXS8yFBz2EqXPffW8wTGWs2/qjKNjsXRO4oCxLBEzwQiEr
deqlPg9AMO4TgypU8iZ7OTAdk42N++et0kYWjsrHI4fX7YVECndzHwNghHOWpAX+SP/GMR9/yWAZ
k4ZO42D6ytvWICMFRQHkfgEk0/qLYcvMsoYHuapZtmXfQhO/2UywW82Cvt9aXSALhGjDEiCSEvJu
1rIBbyf3f3BInT+kd+mVokG5h/NZ2P8sNcpQQdbyBdiuYnaLnfx9eMUVwdYAFehGgXsLj/jyMrgL
TY6OzT6VXJNJpscLZXllH6nQr4JPtlwe6qz6d+xBh4/i+GN2wjdSQpGxIaZ5M7yUH9HOs7zi5TMK
ya4b2PTsmrFzQNLKVFAwu4qijIq9ei8iIQ1JC7t+E/SunVEdE9cWAVkb191hNM2Kq1zZQhsBzQJC
6QZ2evyRcCd6jwCDnkcnoPs+nVhnr54+zAa61aZwjH+tDdqm4VrV0G+Jr7JSsS+qkkk6hW6OrADM
JyY3sVvHAgGhDms6IL0TVMTKODZ+4g7bQdxz+lWCnjvgd37lZzw1bMiDAm2VQ7uqslVgPTQA6rZK
Vgp12/7PlepxBS7IqT+8F3Zb57iiyj1wzGmvz4eQNryTlZwzjdC0WdQtp1OUXeaxPoN9cY3xHW7A
StUfM/tE1Q6ObdSW4NuygZf/5aA2FiLTdRKl2rOK+ugeETi8EqdhJhlTmRwwZjTR7bEJFcZ1JwbL
60XopYAQAxJoSVbyffOm8+yncNvd42Gc12u7dHZsYsvNHRzaOKTLSxybUcN6zXXbPk2U42u4QWQ1
4TR1om7sQPB6fA/rtFlDenVlGp19MWIaOrd4TeaZKoQZfPiiMKWFkJNRZeiaRgYpmIMt57dwgVX8
tdIxdW63TV/Xw5YT/rF14ma1lKRp2C9gwLzQ1DWCgu/FGgclmf5562j3bfu2QCLqlbnva4IGS7gO
p2GpHOsbhgrycUaNSWWdHNqJI/ZqGGOs3k72in35Z5sQT+eiM066ciTmcybfOFMoanNz6rR4zxhh
cRj6yzSiV5L1VR/Qg31s/lt433UqYkfHcgBP6XPBL9zpI9rJY180erc6qxFNHALxSF/kVQhipOAM
YfVB4dXxA3C4sv8ztFs0Sikt1vcguL1nIeKOwyARuL7fXQECVL/0SHcc0+q1EFeZaTxn6yhBrTI7
Cvl7vpMARVZma6GgRu8ol04164TC4mJlnqNB1iUthAMjR4bJ/PiN5JH+8gWbJ4XfJ7jZRQsy7ikV
2zbi4aM22Sezln+8pxTvwQ6pLI2XKgvQTraprKeY/E3r/+N7KOY72ePWs8XNaO6rd4tKQRGiwGRp
KSiaAzlXSDqw+GVC4ku63RQTFeh2tJ/9FXwNsd9Mv4QyPDeGqbBYLok/LB7vXm0hZU14G5eFYG6B
3wB/YJonk96vIod1IPIQDagszBWD22LTSRYwNF4E8te6g3S5ec5c7QJ3BLmZRQgG90U2wRTzcpWL
snFL5CAzo+3elSQb4wkgxnroyClzhB8nxaZTpRQXcLeFA3OZbM5ilPL75ph5FlQH3uZmQGPuUCbr
ghu+c3zfDAce06KNE0TGpWfdQaPYFGO9wUnfCvtrpqDYR+3tYAfYgu85Z+EXccau+W6LbCQOa1y4
dMJDzBctCsMi1wjRiOYOQNP22J+trbObIaVg0RQMer5g+l5WeRqCGWygioY2k8cpbJ4qQ9wcp4Dx
Yoow85T3eiOCRNqtkCR+l405BMSHYQNlKaxPAbcp5sVkuKTzQgtuljUldu3Xxr/48HHi/YcIk7hU
kA87jEEnZmEZc7+QQSZ5Dwmy1bsNsFSVLQ5uc5eQJrDOoPiYI0WyC4mMEP5RH2zGGttF/CWVHcTC
9zHv4Vl1qThUc2tEffTx9MewEV/2EHlg5goAJcqC777w90c4WTRHtoHQaeYFZWzdjQB874UfW10T
kBgPitrlMbo1A2f4jR8tlAZNuoXAIFh4u4QVuEiN5/6f9mTk/G4rrrr0bGv6wRH5XsT5KVUn6jeo
vG0zHFlRCJA/6ErypPzuAi48O4uN6l1ci78aZPR6qLiCVcKQv9Ik+752Kr9upOJAIo/JrinR4Gen
G2ijsLyIIwwZ7xOFQh28r8Zt6PkX4S5FwjB2IooO4P5MBwVexWn5E3aFWFxtV2q43cUnCtaX3n9z
cwG1OrDygwuKWRxHsgagueI3YHh9XwC7Lo+NX+GQOa9k6s9igdFl8ldjOiyjmvuMHNoOO6GXeJkQ
wjFkSN/O6vQeKtISCu3pzz9T6zTRZZV6Geu6nSnETtptf3bfEIPXeCOx5IWoZIp1XKZ2IwL+Udy2
T37NWTWmOdn2w5zg1wfxpWmxltuD+0agX0ke3hy4P9bHLqOpFxqaKUFycxKMpjdGSYcROlJs8VRk
jcA9OtmpRs2w5bjH2OZHuc9WjH4wT7ezoSll8HrZLGCTkAVo6wU/bwo46fD7zACopO2XLrk8SOOg
AuWrljcH4iENOQtXCHuoIDcyAMEw9Ep0TwW8GY7BeCaueH9tDZA+GvnM/9IALU1rK8F00sZvk6Zd
4AoiAtNhS8KtT/A5RWhSINCnAi40Okfz2MEzzrsaVQRvgIvyFUdrknNSclm7J1JOWc+kou4I9Q0X
iQtyoAKG028oZVRL17HXjd3FSGYXxT2waV6iGv1THDvmpCmTqU0S1IdVU63tN/j0hNHHOpXkQJ6R
eEQ5bZtFFfVtCa4U1O9C9wllX7BDpZiDj20BtMsc2t3DvcYKVvWjHX0zIlhcgUwgkyFEWb4f7OcE
tN1XkBmZIQuDUuqootYWOENSxEYOgyGT9dVgZRnlbUi6lrKabNFyZmQBlyujsQG3c54EYwf1eGKo
8V7vOHrTGqdhewZtZNfcicxsvon2Xrtuj7VQbbNhOOGeFjRoTm1iFkP1LBGmOhcQTBtyzZrKYLAp
0OyPQGkODcVnQaFTontFXF6wAzoEvR4iQxY7n3B1aZTANkf14AfmJtU4okFNG24R+5BorkCAF9mC
GLqNadeWHAtuqVjt0gRzubKjaiQyiy7nCSo+FFBZWs++g27cFsekS8F+8XLqZqIt8F8J2lduF8me
jpe+SU2mCY5dtaXNDwNjLxS7LayCFH+5EAq0OgBPbm2PmZrk0CIBME1AIVJO8tO9KDk+we5IF9ff
/JcmlOxPV3Il7Z3Rq51CUf9QS06IBtWDZzsqARwmQrxiE67Tfd+oOhQ4wk4hc4hHz5hC4836JlS/
Esjo+0L4uK5sZqKy2Yh1IHZctdq2dyl12fVDaTcKq5jBMs3+twervbEFb6JUFw8jT+B4lgVyXjw7
usykCj/ln0oOdrP7XBw0twwHTey/dZvkIOrjasrhXBtupSndFHuyllHMTzZR42gBQeovuPCbUb5G
aUPLUCFEjqT53liD07ke8D1mntQILW4ZnsSbatCg43OM/jnYuOl9j+A9apnCy8Hqp9xHXh2O/xK5
jJPNundHR686YhphZzLDg6RrQDhl6SrkHk8f0gMGQmYf/kRndYCkaMgZnntNBgohrdkPkb5ne5HG
7JMH3c0l40AtHST5u0fAW8/8WsfkC4LS+Mh1V67QYThS60x6+ysPTLoLalfMxrrFBOXmZLTIntE8
c8t+bt3oYQD0adGV+aOM7O+IBTSFzPly3W95OQWO+H5o830ftB8jtcqQOZI6rudQtYC6W/KI14+W
7LalgEWsQX+O6qXxsYINs8/mr/jDxoRQzR0VkJqQmjz/KhHOqM/sVnNVmghgxqOVlgPEf2skzw5K
O6stCm5Cy7SS7U5sy4Lw0DyMXgkyi41BKTuHqfI8Gnl9HoyDOA5InvuTBZKcZbzVQ5Z3y7O4I1VZ
P10g+C4rDK8CKuWhYU+7jXonr56+LIqq6gIRdejYBYlwY3+dQBZexAAFcEaiTichNr0eCFHxbUgx
LhcBcF0FU2sHmGjjyDpiIwd4KFZZZhxJLCoT9eA/G13kc5sgGYCcf9ttNbr38O8+nYxAHXzShHDr
iPD8fmXdyW/+Ihu8Hub48lbChRf2O9XDUEXbgMrCY/jlmRMdsLAKvsYns/6RgY74nuM+EWiV1fov
s/OnmJkWAQQJKe3g2P68+8+emq99gLF/kzwHFZWTrdvytAEZ/4XLCmP5YAzDE4vJfGd1+XFpOUgq
pGHoaCYz9f1ofurS28vEAKL6KH2MDBakrjnNI+IzHusVrLgFLw7FJd6neJ6MjRliUsBQkkC/8gvb
zBItmMVaAOTYHVWqLdI+8HCETQ566qCxK/YsrM6PmYQEN088LFEu1YFZT4Puc5x9cws5s/rqNuz3
QnI2UEdbOUdLivPI85LxK2Wmcz4NIZyJG3wj4+773Oj0+cdGS8SC9P7qE7KQYR0t0PrAuuIDx08T
+ybqr2yQ++ZSIWMcAq8aU2N5QtSTmYemr2VKvWUblVas4gO3V4OsjDZLcUZ3bRmLRjM7vIfd9eH3
wt7D1Moas3VQke5WUv5BRqLmdp3qiGhKg6fNSEDjqxfeDPzC5evQAtLYd9aVJzFqGJlCC+8N/LMl
AcGyn10QlfYPZhk/Irc5SxI8JnNklI3SacYUe+T7OSGlSCtPhhiGaFpNAy7H1z5T/F8gK9BLnri+
DEMuKcGbTjrWsxivVMEo4L18zINbBV9ayHbypwfP9VYcwzO7SNz2GGx3jU70IBDTHdN5xoM/JQCi
YdU6uK8gjwKAxwQVgBLmQ/PguBRDf7QSOQUtCpYfSierYQ13WOYFnmIpQvdkmLj7tJ9g2gulZEXR
Nnd/S25q4uxByIMR6wIXG1rNM7z9SVNRkK0UIp8DApRU7AvF+TpRlgXr09SR7tIwF7T4sdXQuaHD
fvZ7t3HkR4jPnZBP2py94N7l6oNSrPZxKWY+6UNnuX+7NVXesF7zkIY3OxRGhNLO599LVusaCzYU
WcfQIjg/ljYHxpToj3hwjVw5esaBoDu0RZgg88mX27c8w8dxKGbUOpEylldHnqELTLR/lPCTGMcY
BIIcqh7BZOlp+oXd7obPF1PSK6Be1xXrvslw37/Xfva4GVgZpAwgR2uUpEkqpQ5IrJ+bo/E10Bmw
z8Iu9ujXyWlguOLNKbJ3O6tFUHa2jNTK8zexokS0AxkdBiWW8Pr9ANS1Prc924ElIfNsVWXEgCQR
050mCRbcxcbodRsDqRIf8Q0DAKkMUY/hkiOyAhEGDXq86l4//DthDeVILsLU+hrcE5YRPn9mllpT
/gGujqV5SgL/2jw0kygIdE6cR/dgRzL/YySVZ8/XnMsKnI9RHfgznvVXP2AymfzHJkh2TypPNrDp
oqwn6VeaQxW3+G+sj9LuXBI/EsIOmH0/ljL8NHH6MLvkjnPu4Q5esTTdmBYriKWnjK1QegVb7W7s
Z4St4PQReFrjaKitiimfPc4h30680FRqhQe43zw3j/2cnbdnjkXQdng5BSJ+/h31ZOUPkn0oDztd
Vus92Nf40lO6Gp9KYJ2aHpPgqEhPgVizMZQnb5lJU/XWlcoaIYSR0xPrKlxmIjiVinnKMVIKoXZR
YxbhsnwzzVzidwNcPcvPgCTrcTuocbA/VpgqWFbwLEElDZS2HHxuB274gFjqD3/z3syAUVqgmgrA
jc60M9R0CppS2fTxLxKmBSinyu3SDVsB87NXeDTSg+bfpi/sUHcAOPRdzsjEbOhIFqwJdtypz2fZ
xBKZ/pP6ejEdvhE6ynEW98lITreKfDiRdWAqUpcw7ff34lJ0JAGdjr4parWqKP96Pp2FprsKNcmQ
3rG/c9TOCfWcTiI32uKi6d9hZe2DtPmLI7k11GItdEeerqXUNZXfcE5lSUiop4txeh2QnGjEcVqD
/3gliNmTOsrhUBad3yJ++F0AsjVSwRtAQgZkdIk6Ed8qkLn2nUFht2UYYaDy4rOMjsCXUg3UcdYH
AQQG1YlMpJmr4qqfS8JTYHxcUuc0ThA5vegQ+vmEVS2Mqi//DJZAV2/zWG63MIi9B8ENB1UIqqFE
Ui6loq+4odw/EHM9gGSQfoeB1I1eP8+Ns21KEem2H2KbP0NKSCfav8Vxn2F9ov0j8OqPHPV15t4V
uvoxaXQZX1dM7/5pRwnvr58k12PzpuJbggO8JYktAfrdbyCNqFGcG1m+/PPyvUbei5ucB0GkqNZQ
VwV6kEe37NnnmsverTEvgwVlLtNyBQqcMPrOJTpRG+yuPwv1GkFX3wF9NuT+cV2/Kw2eY5cIY3kh
5b47kGKNqtdUMLDSmfUraUqiTp7pZ2F4O0FKPddNNG4KYi6/wWsBhC9gzjQlrqgHwnR5qZTRvGXb
/06/O/VA2sV9rxdSCI9uQqFy+OlNSsyAMRqpsP92HS4m2/9Dy53/vsTyIeopLT/m3ZnCH5v0AtoZ
OatiFPSs6nma8WVlDKVtLej4+CTktSrl7oevoabWPmUuYVsCh4xw4DKm6QLyhYGcWj6kCMEAORg6
mOnM4YhpIxbPGhpj6xoBiuVZTaVCyvA10y5V73/PxWS9KfwjtkT95CVZlQv89P5dfPhZui4fhtxN
Et98qdS5xntRF/zwJdd/9Zrnu+4sKqK5qV4Owr95FnkdtzFpW2xgW+9XRv//OF7LWr5agLMgSkZG
QLgYzxNFwZmnbaUVz20HQFxamdcvUuEGyd+EgSh+QaFhnuAh11zrzTx9TxtrXxs6E2LguhlRpDOK
arcEfjGlIG00nTsmQ3/NgZT+tg4wxXZxripU3kYjqxTpMDNk20NSuN+/pes3BKtmQ8aYlrw3434B
KXTT4ZR8FbZnJpYGzio8tmQkXBcp1Gg/UIezPCOeq28ac5ln+0aKAd2fMzDHkoBL+XXBcmLrpzDk
4AUe9WhxI/XpoUe0OZai3dG6hgcEmap4+k3rYi6koUXcmprLzhN4EIXAHn6BKCyry0V35U0LB7gj
0k6J9tm5YbAHQ2zMxb+FHJoaLZVbpCDixVjR5uv/PnFLjv62Y0LDo5Hychn9xXoVp5NqYYyN3PXv
cY4ykwb2QrahQnDUKCuWhRKiRLESQkYEvf6D0v0BLrvF8gIckbaqHjirEmk/qJ/YuD7jIKC13uNg
STZNkfdiSwXcZ2Gw6kOUAV7lHex9BMV5P2CDZPwH/MAwz4J3pYGq9I/+Dl/iDCUXd/6h0j9ofzrw
KTcMN19jysArQkCIjGGxUlRZKPA4DrF5Qf30kDdcKgMN2QgaYrass/U21gusu0Ndq6/hKPZqufNF
aCMK7Wk5Iy7vp9XymS9Ph77xZAP877wRHX8aIt0VzWVqa+MQzStudnGPU9TCXZFcf4wJC0e2OoNR
g54YcPa9OD1sqINknslkmb2aOSnptwm01WJ9p6vRT5ktq3GV9sfj8Fv1Zy2+mPAzdqzAprMxnXlZ
vdfjKPQxt9ICMD0L7gOLlhBoB8xXar/SqDQ+a7NZfxmyf8Y2i7U8Gict8OKCRr3arlxRaave9fPh
RoRUwzEPENE05FHnlFO2MxBB4G4q5rjru92xHsOX/v5Qw0eahiIxZuVxGot8A3k3YvSwuvAf9smU
YFSYsQIdBekJJ4ZKK0Rctyn0vQWm990Kw7kTPDSva3FzkdrhGMqHVtltc7i7ciJNiXyPcsbC0c/l
gQNSgggpNgQhcEDLWZQdDh+0PzIVFheSq6Gck1f0rS+1Nfb3mQ0KfCpODEds2MqhLkqH0T0Dg/F+
/1FqfsDwrP/vx20vRirOTra76SHpwNeprmbpbyIDqbbzS44LlKGWYzYVldU1ssBsIc8dY/biHyXi
/LnyJQe/fmTOmFWBq0cdzaj0RBGa6lyUpVfb6HGt1xEr69utS/PILYXDlPPvG1k9tvgYNxnwPJxP
s8+yBTIqpx0msR2IIWoOdTEbHn1zcx3E6RXSehG79/XdA0Ffi1WQtyvXpBIOTPBFsnWFmwgDI3kb
8MAZ8CJ7iDdMcby1ji7lEznzvtpFjsJGClM47hnPGRxLdiC1DvlhXz+1qb3MkfIcOWcCg1MfuttG
Po48x0d0Mm4/IOQdnPN/Yyms62E1TeD1BCxmTNOHFjVWB0y4bk7alLomthGbVFFf/V6jB8ookaHI
HSCUcwbLZ3akLXQpmABsMQ6uQhRbqtOZhPhOSQvdS9KB7+6IlXzZKGuOmEqtwW7El7SGXNfNxxHQ
cau0sWqWCBiur9IR/jZSLgGS2dxLhz38zm12koiyKLbdXzn8G+WdnfGAHtrU/uW86RNEH6WYsbo1
ZuRlqzPJHWUh5exsqmOf4guCvnEVRFfvIZt6YQxln7zPafBLsFvW5KNaGHJ2yqomCH5GeVaix56/
yHyN0b+P5y71nuoK3I9CrR0w5aUTBoFNHnnOemqKqglkSRp1JMx/lbkY2JUPHVsWkEPCCpDAfypt
cPUTTgp9R+9PRorfMxOIOpRLXXLFBIZEUzw7wjYToBO3H4ldeAHjXXyGMspspCKwzqmo5zQiGDwz
qa7nIwh4OCGYPu5SCA+wkhB3aTktLa5OMnRKHlMb0Wjb83UlYtMsLI34e3ur63VSseTd1WrZNKJs
L4FYSmfDzIGSwhhvcJeOj9Vq/GMJOcPgpP/CsppAx/yNi0sxFVw49JgJoE5WIOgFAAHOtx7y5hV4
mTV4GuYxq9875e9ZEnGBemUs6FpLuP4fQa+HKa5QSs54NGW1j4X/81waR5uuT7ccoHGlLROCBM9A
ps/UrylZbomKZ34/N3hCNTHZeoAITf7EGXcwQKbSF37/CLZnEGDZ6wH+LpYuP4ZMaHVQCcIZsSql
w3WQGLq77aPj/w5Qv8CPiutTfKZk46ATtB/w7bFTDBsfmm39PVaQwiVIgyyfxNJkj/BMPqd5tLPh
OQYZpGbzbIv7LNfHMtBgzPlvGaEMl81J4zGWt012/EKL14e0syzU6472YgVddfBD0NTvFpRlNYLf
bflFX3y6qemFPjBhmE3XUuJiDkP0pC5bSxUIbDer2RVrBvARPf3R2Jx4BPixscX4kQnhx+ZLw/RJ
d0b98VajToynyRo1SQq+sxl1F1V0wP0CT8TNA99piMzwVj3A46FR38++IiI3smEJ3Af+QkyXmeLm
0DHsbjv1u2Do1mdlea6WG1OM7jfPFx+KO14Ezyo9ZN/Xuoyog6N75AXKv/23azhCPere/pSbmkSd
YbjN9fFz7Ovh1ov14OoDzNyeIzoYZq5nxpdRRdRNc/1L4ssiTC2yGzKkTvi36Ze2FSsOJiS2H78i
7alsHJ5re6DF0wgM0pO0mgoKuR9EuAfBTS5tIz7yYbAGTlcVj5vJ73vY9Tz6rRbQQ0+2peOvoIIV
2eBjQVG/Z0JkC3qEsRq2FPEfJz4+27TgJvgsLozISgAI/q99HNQ9L1tdntjUOV3xX4ToxV0IkLGz
Qm6mTrNGtjwxrPC+6Clz0NQ15PgDIZybUFgxMZPWjRPrjQveXOiOqUAslRhXsoxUIQzIthwU9hqA
2Jqus0WPpq8AeyqthhItEmN2xotfEGr56lG3mmLss/OJWV+icGXqn29RI+v3VRM117YQrmWN3iZu
OIxfXwU7f1grGJ9f58HqCcYiv4Z4yWuSM+Wt/H/MMjojqjRyssFIpao3zQi4aaJVAoB3x818RLfg
Kuw96kQiGZnZPp6BMemuadNGovW+FKrbFYnOwZbBZ6beCyVgVx0sJd+KZknQxdd6CWUc0fCsfl/X
XZdDahJtatcialxMGaezyBOWu1moUD5w++HkQiDVNbpCjA3BT8R3x5AhJQYVLTADnuZF0T5CDj3e
eJ76Bf7w+2H5jGIKMnK6lwd0g4WIYDYEchFnPppLwuAoWhlFPqm+o8EIUgdHvZDSZeCzgcq4gZqU
shWg4yankVxlVK1R6klyGmH6nyVVfY7VBrqCm0QnuwIYYghnQA3LJ+gboJvAcrKC0iVC4Le+emux
Ztnah7Uywbcwr2XIOv76N7PgTgnahHJqNh9kPbYSBT2vARpyRMP20VA+Z8EAEXiO3Pge/MLOClqK
PCTNSbg6iqks4OF/bfsOGSHDKEXCcaF5t4h2imdZmmBQnMRhf4gWgEJ6LPYrJ2s70RvwRpJXyFVE
CoQLfbtSdUtyZoYcXORw5t7UJ78Ke1peKc0sbv/EltnsF3t9SO3+7227Q66xjv4kh22tRODMaG33
LDkRNsqcvOaap/XL/h7GpnQhcpWUMoaksbK06eZav5kiNeUX29qGycmR7ugdamNbrERx8wtnpb7i
77gHP5GlLobKPxZ3N85uVS+qIPNS9TKkVXNToUJ5WiS7yc+cdIbCe4jDiZAehZgkDTPHV93KCjJR
RZCl1gVMaWm3/8S/KMyFp5fPiPImvMSO4B4qFDvb2B+0QmQy+TNZTNPEIyDUBRk/00JwMOcrcBlk
+ux2Xsf1Cdgd5vIdtoyuX4sQaFrKD6myAqIVlq7tV3lAgJjA+G4WgkqfssMI+8z6uP1c/kzKwqzd
dwCqsQ9K2iXIK7c0qSxL2Gl1u+GfF9F9AcfPZn30eJ5YzD3YJ74Z4BZSohrSkweqyTtBt7FMu8z/
nHGOl9kYKcCCQstZILve40mzXwwuItJng3kWaCoyGJGOWR+K+s3dalGQy2ccKkEcoCwf88prPDLm
H0+oGcBWGo88sR63IWTkVR91Ql1dPEyAAlpvkpjBrVOSqcpu6KKc/7/3+3V2ZjRkXP/Bm9lMsWPe
ydq2gaJvS/peY/kPF9YGUcOSkfKE1B3hiiT+tef/9Ceshk9RMCJ6Lds2pfRVxZMfRr+6PvwusQAi
WmPAPcT9EfGgM6fP5Cg5rmeE2Gn3iG/yFRWi6WjN5TDXVBjR0qD3WkygFO/eo6EElRqOhGvESier
g73zcLTYzEhFyAJKjoGG2qvPZyAOiUfvlGhvyXO9q2qcu9Q+FOaXOMjw6NlXZ2umPEySfWQ9egYs
bJ7rLK2/DbAPe6sTcEArC86+eEe71cBSVVUSnge/cnF5TZXJnyCbfdkBc2Mdd/Emq5Zrgz5V48XF
o4E2HNaNP24GgqXUKxlcO74MfRT6Bk6Y6ylcmCOIQmLNGpMfNAmqGnIVzr/sDeuRQ+Q9wu1w0Gck
g2wNJ3+z5HnwaFxlj42rkDsLwRbt5VOD9SpUxRjxqCVc7vuIRUx8rqThkcWfb+nSy8AAE4BP00eT
OgjoSJVIGOm3NPvy5K+YCy9vZz7OEjs1AlroN+AmT+Z50yCskCmM/7DVzne9Cif+UzGQvmcsBnIL
xwWFdRnk19rcZpfZ1YgrJpW3zN2rQIOwUvUeQrFV6QQdMmmuLD0cjVYAkCoqSF4njJ5v9j/zVKir
5jvteWWGsLgUIdDcEGwIPJ0JIhy1lb6rypAkOiNCR8V99VSILAD037ukGUiclnMK4pMcIXsiLhCR
cntjIL/cj9/whWaN9aCp6+ZzMcaD7i7bbeuO7cFWMH1zpzhqT9/SKbIsB2jzN81BpODCCtgrPE0x
Iwts0dvRcyKZutIiCSy/HZeTz0HboTVQ9ecuP8LdjMELg8T8DiBo3hygtk2qeKoSiJiOf/7mRlUl
czUOciTa+PHdRZDQO1yU2pVUNJdD3kJg6yNV6PTfU8k4ESDiZ/m8tzk7n4Inc6Mx3AX6eBPnlOC6
lMh4Nf8fV5FLpy0R1pPtZYF8uGnR6pcX62Hu5ttoQryZv7FVDxy/QezuXD00/0S4PBseA2HaCjCy
XYFiEX9R4pQe3uCgtrZXgwoBa8cps78MfkwWeObVx3QfBoGH/H8vinp88D0hWg7ZDjUFJJyiK6Px
eF49ivM9nhIUDLFbHFg8rbPurK9x8O1IPObq9adPQQf7ufvSeWG6fj/DvNE12sr3BtPxGufoCWIB
KIcIZo9Ls8wson8H5aY2MAxXnIx2pg3iE3R+P4/dPxb91EiYZjn6LOEeYVBOaKG7Npe8Hwyil8VP
gzOtWqIV6mQcDo43uP+IUXSJxxgoCiwpNXuW26Mb78+Wo6t5TTRyqcxux0KpfikmrBm9MdyzkWd5
lsuJwAHsIYt0p+5Tx6C2GPk1y2HTDYJHKgfCgAog+hoGXzZhfizt7sZx3xXeea+hlN6kdWKXE72K
JxCEgPeGfOYXrdGNkzL4zrMp+KtJ13pPF/XZFvEde9VgoLBURdnivQ2xS/sluMJRK/aV9yin1YKs
t31lDH4zccXIv+7s6X9ixJbeCCpwgUZfwc/2/RZzCTeBCBJP3Fi+9DNJ4yAF0791Y2a6dfl/0+77
5nYQoBmlW99ShlR71ouFpwhPr9oP7EeD5T2T7rBseAcSAef7nDroc89fj63Nc/Gs3huRzOeD7KhO
17M8erS3SQeCc7uV3c0VjAt6QCJECaUGe/GRD1RAq3/jW4bEVWGSa+WDpljvo2sdwmKlZKP0B7vi
LYzWbQ/HhiqR6DVdY16PjGZTCIQmSEeh8J9a9Nv1JdIwd6yYGz7xirrykKYFrB8wcnEJXvqofO5d
KVI3c766ToZC8jEAhF/lxwPKdiKZbuqUWIBzKhuyQ6qbuw/8gnI48eICazLvm3Xi54e3mG+sggkN
bcn/MUWvjOZTyUuWaDvZQ4QDUNwabvwm4745Z4XORT+wZlhgugBDXiB/A6vVozsln2iuq32Sgmpx
RMUxEr/IHmyq0Wbdg6Wht+cf0r1vcyvC+QHRhOLhuyX7pSRnbsMMuNQ79cFOifn0zk79QEr39eps
Q4BAt6XvMx52BbHypwMwt6tb5Y+Z7IbBbfDi0ow+0YV8mmXIq6jb0rPwt0K0rOc5poITSQv7kJXt
EhoCf+/0WAuu6AEUrT62KQB3Ou1+mqxAnvmesOoTsFBZ6ShcnzO3JZayOYxsyeCfwhCm9nNkM+58
j/BGOoDf3XJvpE4RJF41iWk0K7Vy6IYlFo/xz+TqEY+kXPTyHHPna1Mb7P8VwTLtCwIr1tdJhpZb
Jp25YVP2zoh7+MFUvQm18TNhWErpIHkZ9mHnJ63w//hk8GUckF1ekhoUqeroSCkL1dTAmYvs4BpW
skMku3UiEr5S49s+ouISm6g3wQTGHqIKCKpQHU8YZsnhHujqS3ZO/7m6QJ0W1Yj+dmBnjgEPePAv
38LRhkkHSrR+o46VNt3GVgcXVO+ccbkq6KLyyDaw7I8kCwSZZi5mqgFQTkgtHiMLCLpe9J11XxKG
YA7pu0SQFoQF9yZK7M9xzo8iBwsaIn8RL0eiYwxSpZCp4s6NIaCt7ulMMzhlKbIwfJx0f4KSrupY
XHWbT2yzZViANb0RRLo7Aaoj8b8GHwOVOuXr0EY+N01+Yj+bZhKhw79IxKTscJ30O1g7DstU28t2
sCB4NOi0m/X5zOlISOyD6GC6X5iiPxxVp07r+72KRqafFG0zQjNLP8L/qIPsW65obRaXUIn7lO2m
qTrcZUD0QJSLuu5JEadXz9ey1Tz4Wf87aRyjYQ0C146pvMZpi4QqkvL5ZRvZxNNSR+f5fMlfi0t7
g9zRPTMYsadBdyNhCmrv4DDYJP4sbLTPZrPOcfqBY0N0NRS/XI3t2HFuY4GrX51QKvO8sQek0jaM
rqMFdI0EDeUg709Gs9tb8EmRVbFLvv1A2vTyKxJ6DMC+HNL+gRyFBe/P4DgeSCZnaBA/wUBHrGb+
VRvUWxSYfxEFOdqWWE4NE3+zbD79wkdlVI1YYldTg16xmtDENO+a5Az+Zcci38ekM9NNeC2wba7G
TG1t97eacAvHcr+3tLDDCaElQKRzprH+ZVh6qK/SMA26NYDmXGU098rL2mI9lxk4nUsxelyPOcV0
jP/EOiechdULjaSMy26KW8lpIYIQp6cXDzN6fTWOsOom7CCghANNtJEdBbmeaI5r/JKIOrheLlfd
5kLcM6FlUsiSPSBaG2KvhtcIO0H21CzC6Ms718hAS+LBDxwZyqDdyWUw4c7fvk1EyWLuFLImiiq/
9S3F6Gr5HNylYa070FScqXjU3tTFHUoYg8ZsC0XFndkb1Xb2fkCBi80Wbk5IQiv94OoBY8wsx8P3
R1LhRIBM5MJG5lY4kvOeckNZLpEhyahtPilQJUyll5w5wYY8rkHQQgX+2a/Bg2SWxJ37wdzsKKng
PoJ5UNqf4ozXe1pGNsedOmSBqw0CycLQGYxopDhI2S41E2Ik/jRTsdiP+BjGEQsxcA0PEjM5/V6K
QgIlLcN+3jGeiPoMR5RE7yXSEXg4xEUKt7a1Bv3hMJ95v04BJqQ5vBwMZ5OubmjjsFntTwbYk4PV
HQqwfE/1eVn6ZdVpu+KvdSEhZesgcPQ5ajXr4NhcmP1+q0vAfwjGvvhQHj7dGiODXIz89EL9xAkD
m2+HO4xl9mtkRfbiTNw3cly9edXyHTOLU6Mvf/ElSvx67otNt3g7HizX+gvRTMfLbm4/shhL8I87
MH2o6u5QQJGN85YqfECuxOpyV3tmUcRaELqX776Yiy1S04JEUXyz9XbhbWTG4UxyDrmqYjSZTiF0
g1ohesh5/QLfU5f8hIJSWTVy5/Np6XDSEPKukb8ZH1VwLIkLUVUjswdEihzSJPyGzVFYw9meI06k
CBcnTjpYlylfuek+XzzdBtByarFxNuHVapih0c2yXuB8jD19QfrFxASHV0wTnb+fDBv3QaXQe7nh
f3GLmOC0Au7mu7PHwdOaxnbI1a2zC4OnGVslklG+ndpBz2W4blWL10u2X1mz99Y6+W145bEjaRKo
MhPoeHti7p0QW2B14tRLzPaTcej9ghK4d5MfHFks82xqXzgv5Vnry6/UqM07gSQPtNFzb1Hv4qRE
0gegiHaem9LtzzVnfbXbQwL9i7IPLQzHFhiGpAWaYSmfFYx8WPcrUY3srvsJwpJGu4y9bUQXum5g
Cks4AHjPgfc0e7zK13viAQTg32XYTj61KmWWc2GLWrkSbKjEZScg75NT3KKz0OQBt3x0CFEoJg4K
JeDGS4ptEelh1Oyqh+JHQhzKbHVFELZYzwGzbl/lzBRlwkd3Gu7QDoJSA909qfOziPmOM28PFTTN
hdqayKu+HdCXeQGd5nnmRfjYXzdC9QHOFNho302DRxinR72HAOZiTzI9/6nUaYz2VcpLvLUDHIxI
JyuSXgBdwUTTh5SjyGr0e+vIRdV25T5npD6ipbptfOHyHteeChhgiKvhGripNAe1eS1FDHBHC/Mu
vPYYHZTbplNCGmLHHwZdj14es7E+rsdJ2FWTVI/O6UzkdNi6ghiSF/KH8QkwPXou6YEQSobERlGn
S2QnI31SvWEatMr1z2TJE9AgJxz4PPbQd+AceV7UE9qw5gbqzZBK9RQ8COKKgfL5u2yNDrkdqgCz
C7zXMs5x09bKEv5zOiivne7xSctSJ6VyrgdlgHHATzg+UpnS7lDA+tcbuE/7UT05m7n1vTJxxFU8
yKkGZ0neuwKxCZDHtrg8OF1bqzrIpMBg6tDaHwbw3G25AABtV55Z0JVhocxZfWuXW50JdtpYYHSS
xKD/t2a1xznKJwEgRK/1kpA3M9VQxNXcneOfG44ECLEtzCOaefINrhOLY+4wNtPjAqFJnY8vgEm/
AITUtexqzRxniV+5/TImoWdghmXT7S7EA6+J46LT2CrWnUuLHiRYL3uomQvgQDtY79TBGhI1Lcvg
yT3qNvjQngUSB6sDRLh/gljLFvKjxJd7X6tDTbOz4yZZ84DV3V5GF0woLAPoATw8tIbkqjLtZhwc
e/RfJuxWfIS61tg0z+I/UMIUPaVKbpyPUcmaK3YgviKe5Sr3XF24YASkdiEfBUjBP8WUQ9i5xRKM
mK90N+IeBkDqBgtG788xpNgUadlXS7mpUeNnAoxfSPpwhtLyscAKox2EAMknjIo25AH4m61am4qa
SiqhWqQ4Vl2kblHc8RH7Nh3vO1MSDCy//GKFtrSkk2j+fCtEukYl2tIYB4S6KjxgmsgRGYsJsAq2
1rBBphzDahzRv7v7bpbGQkQLZzyd0Y7RDrZpQA2Cassg4KPxj5nZyfBFDp4NZYgDahPcIe+snHLy
BQ8w+EA+/GIa+CMV5zyHsUjHg9N7S2sNYXyrbkrvEqvgnDHEzB5Rat7CYpzt+kLGy1muKAztSQ5T
oJyDPG9PStqlWiXY9Lx86kJh2ktzBjOYtxv7Idk5a1F3o2qkRk1LLY+jFnynyhQ0/AutLmy2Zq7t
g+9YYu18U3VABOkGYdpZH4renC71oQyJ6GwJqb/P/Va5cUuu31Lk0/e9bbGJWQpKPo07hgL1IE0F
D622F6b3JP31jcVpPlN869NaPVonuPW7TQKf4IP35Y0zK3BXyMhROjdpAKGWF3LdWbr32NB1AOtu
OHnBtVTmj+If9V8rUsFNnPzieM/fyw1nx4kirBCRWECcmCJowGP21+2k04D8iANkXRZ+bkxaZpKI
KlhympXFUVPI/0RQGK5dSQGVTtPbM3vkaTcuY36QEoxSG/8RXp4ErqnxzvS0aHDKbMrGNAPOgLHZ
cSd43xk8z4Pgxw5InbsLPbHTAg7V4WJfpZD+Q4X26XyPTu00K+JCBGneIMAV6Uh+/LRNSxenpeSl
+ELG+9PykleTjDu7DzI4QNVOGvO9Q4b5TJ8OPc490gqly7H3zBSXirOLXkYVjXUrWuKRRhnItVaU
sEngLLNQYa5RMSpNwuOcPx+sGhPGUd4DpJQxD72/pFgyv70h7ZAtiJ2j43y85lrZxsnugGT0UROf
Y7I28div/p5QOgVGwgGBOUUiMP0Hy4rZY9cri40j4DS+Cdqma4bTanR8Ii/78VOqDYel4DQqGuN1
YgbdRv3Hxfr9uRTRo0Y1Am3mquS9AzO4rLlxFeLiooNFjUNH/uBJic0EExtamR73p1CTtQa5nlyz
oBBxaLDPNucmj19zkk7oEB6fteTqzvrG9prXysHudjdF7Ec/EyNVbmDkgO+Qx5/042MPi1w7OqAf
U1fGD+GBOqnvzLhp8f2TjHPMXb5GyxJIPskWGTrW7rfHSsCJMEzyDCnd5KlJkANyS7XRrhdqMNTB
guvPVZ5FqBSEnIAdpTxi79+7y4zTFpp/fGKLpouBC36pdT7bwDuT9K9h8IbKAnilAed7kd4AT4Yj
92+QGDIdr+lAHmpsffcEtrfyxuBEMhL3fX11O9V94oMqPyMkLmSH+aeSZTXBMDf7objPQvgwyvsp
9lEyN5CjyWVGWSdlHlJx0svxVIf2hRLFmMPJR2lbdjbajqXVq/KIbk38VtlHYReiK5zQ+J6rye8Y
8GYHtOOm6IjN5isrn1VgBP26qLBXL+Da/UhPYnbiFGOtolv1LsxY+4LYzbgCmbnbmEbfg6TsSyVQ
OR703o2dak9Xo73fZHDQZLZ+xQ+ozNp1m80/MKr/LeZXl1xhTYVw0h7CcO5MfvwgDm0Nmq9p3rXT
9mSXAOcOS8Yf0HowvXOMwKFCv51PjEnuh4iFqRCpIM4hhuirUQ9qAStQvOdRV6bOjW5OeqVTgZOk
JwkLhBGxynSapZVuBJHjvbtt24eg/9wQn+5izJ1MXfhI6Gvzuk2IwbR8ThPFUD8gX3u8uFIBb8Ub
tbM+pL0bpmso8GQEiwOW9jzBV5r8QHFEreRcw5hkFMsQ7Xi61GumyVO0FqjAY66ViQCwKgmsoccC
C0UEnof78ocmd1bXjNcDoM49jqkD8KJVN9IDfGki1S1iJWvScbLYOhS36/qvUWGXXC8e5RraGlzt
S8uRAeaM2Qh8QX34if0I2xT62N3Iom1QOgTUmgyW0I3SuvvsA5HAt2dO0ErNpCfr5JRA6F94osQl
dsBz4ccMdiPvZuH2u9DMProZsYEPFqr396bYEyqvbK69SeYL9GHDIzTwVg2Hog2m7LAmCGRLhuW8
5iUUv+3Ec4/nztZDnvuFk2QTXku+0+NeMEGBNMGmwHM+nzlpiWH6SQJlToymORvF91zfMTtxXZ93
RcLoo7UWa0pVlg1revIKUkcNUcrkWY7n+bFO7PFf56sr2tNwqVP5FpwMC8Il/kmY5nJs42Br5s53
SlTDo9c66YRY5Yi5N4hm511nSyG1PfuI+f0NbrDjhr3j12eNxjqXH2tUnRsJxf/ctNk7p29oo+1m
CUNHNWrSfeyOUAv58J51OwnYIB0vHvghd8vozALfm8RE3+Ph0QzdChEuZcJtWYO1Ces0B3UE18od
ArTyEKvtHmO24cxbnNUtk5w+Beg8LVjrTvzGdGPFm9+jEteMGmZf5DtIeMQeL4WSjPV6cyc2jSM4
F4jdvbsN0OmgqVa+PsO8xA//gFomUgF6IRFN2b0RCLowu6qNkoTPOQko5sg6w0PJUSWLJs9P9t4F
FdyflfT8noUtxKYI/8Ok0D+RKaRJnhtlkQVCbEQb0PGhysY8zKCcJ8PiyybTxvUOitLJ6xzx0JjQ
lMZ5xQ8qhQro5Y3byC5mUeisPOPO4Y3InoiALfftMWYGrwKfhx5ltRZIKyNHT+eva//oUih70Z14
KdSdzQnA2DG7peJyevsk52xa8e94QV3qJm2qjytKdb/R6LPIPWEewstkwKFht28/n+G0a3W5x21t
YndsaapeyDj3vOkXJS/y/HvdFJysJvshTSDaREjYriSk7O5l1lHOIli3u+7ogRBOQmP3gpQZPk0S
Tr8GwQTj2m9WQfGPEb4UY5K4PYIpq80JVegN7OFRWoxJ2WeVSI6S5iv8Wuk9QB77+VkAlbRl/lP6
NqZhHkZ5w9rI+e5lpex7AwPafh/7j2jPYAzwENuVhnr9NKy6ZgsrG11na7kusl6+MgV462uqQbKI
5HRxQAHfuKA9AuBef/jn4m/8cWT3Cv1KJ9RNocZZGx9mKr10cQvS/QI/od9o6hyY0P80y5I90LwU
8DdqERkhXfu3MXH8xwVjJew666Kb8Zo6ZBe7yo/4ax91jD0B0rcSrP7SK8X2PI8SR8OcHU/kdBBX
AmEBKot9GPr5YZ1OjPCOcumwq8RC+hy90QzlcH+KcX9/aR83IawcVkEhVpJlnhQ4c4QVulXVIzra
0v+voV4+dmxh+G2tKHIe9nfekCiINsNcxUqvQQjC73JcPoiocaA5tkbCyNdUxBoTDkUavuQlWXH9
dmZ4a7Qt5lTNEypjvi4iW15ssHU7dVThkFW6+jUtYSARaNnCuhayxiVFxx527i3hjL5CkLDZw0wv
RGc0vfQf3Z3koy4igvDtLpTIW2H+0y8yt2ZDLACxobgAYyfBsWUf/EzqwQ8mo5F6rmSYl03wgkYI
TrLg9bwr+V1MQL02MzyIEQXxWE+fvZctKlIKcLoo90iaxDT3WobC8DrlkaspuLt4cZynCZ6CBYRY
zEpzsWQ96CVXywk+rB6XWJhfD81LQZK8zJoV6Q2h5//5ZurNm5Mrq4xVM6LuVbc0r9CivMk7/X3U
641Bwv9hIGB7mTjrMWGfbR9aNe/V/5lpX6R07aciard6ID9roXkTOcwfaZrRJFIGEhEiEH0Dl2r5
BwqWza7bWlO0+Z53OKDonI1tK39rgxQsgMs9aL8pNMhtGr2tYmJHqGGrmrP6PDFLAyLs76wXFdVl
V7a2m97M6V9Twe9ZPfGuiOyY3798/zo7IBSiZgvC9UZsOIQ2uM+uz6jJTHZ4EFDlLNy3uQfSaAV2
XupS7veADzg8pk0or+3P43CJyqu1uZ2q+X1JFSIezS1sM///G44nt9RQEbo8eQEcu3Q82rj+ykZq
DckAZG1Uwfrb3cZa3CxLAzS1R5+9/Jimenv5ObldEJkl0D6FlPKRCmhSPB5R+apVLQ/n4vIsByH2
o7/Rdzs6EVKfO1qnd4pYzkewnmsq9id9ii/vZ8T9Yldielw6FVO+fv9uzuUy+jQ25jPQNBrqaYPI
KODXwRt+1H4GvE43VS2HcSUKYmSRMPACVkziQ5/7sgXwq6oiXY2l0kE6RGHZFMuQCWTqM3PKV1iY
dJz3Ihb50mosTqlnXke7+G1qdQImzPebJzhnCuw5831/1vlkIjxt4F/tbX3jb4+IiDioD/v52G8q
wPXP06NRgJNzIxLKGWe33x+3o8Z9eTyy0Sxog1Y6AWNIhWRosNcBkxzNHuglFJRVsAXjMLvNb7Pr
BLnp2neea0e4/LPMKWqkz1f/okZ/mBCViiyIUz8z9jhn2/2StbFNjIXMTrsgUUsnb9boBbOiNwJV
v1EGTQUiYRfi1IqN3c7dt6DngjJIrRb303yBaoRLSbjxol6Tk6YoZGVNoglRA4QmKczj5PZQylzt
al8hjYpHgnDP23tqMNjQjxT/L59dqHCSj5QxVNoebGWe2tqiUwwdCcMpN2bJUgTbC5SRnPjjGTBz
Cuf1Y4yySgE8koJSzmAyiQyO79/DeMq7LM6EzCDWjzooIiwcOpOqAwqDLKhhFeSmSZUB+MHCvgjw
1v2ucMOs/a8fu+Y8gp5HtDR7QrAFIiCTfl/poC44UMU3RfW0C6yRMLHd2JxNX9KOX98u7FbAL9/b
dftV+qD5Ngx4rFHWqUink2KCu6nxILOcvtoIurWKGsZUBY6S1eJpix3Hnmim/Zvk4CyCvUbigkCh
aGgEVfLfF6LVfz2wlxqLUj+1bVolVjGp+vwYwpZ9LzLfrPf+SFJAayHXifaHBDB0Bfd2fQbyj/LO
cDZkErvvEYiUQ/9W2hpmrCVNyHqVFfpNbfs7K2M/t718SAj6SD9m+t5bVfRkYCr1C34/aDWoo/3t
H50uz0FvqzKUQ4cHKVHmeKmFAyC9DNDkymPa5aThZACew5mep9GD1qXwBIT2dOt9GxN7RbyUjkog
DLUYpt1ONzmiMHnRaQpQJkSRW4Oj8C8Ds5QDKri2FsYgeA+R/LAn1PlIQL3xCmtd52cAa1/KbqPQ
NKsUHj+6T75X1lzEx0DWoR+tY7utiWsZjtg5l9EmvDh+1Cq3PMkLm6Cs6ZV4ku/ECuEA/CDYuQkv
5w8W7PdPwp8OANQB/rpXmDwDm67/Gq1Wr+T9o9rhHmW3P3M4j1A7gfSe3ohpIjU5iVxzh3euNhlP
T83kyOwl2OMMqefkQuba8aEW7pqJgKf2OTYHy1W7NpvIQIL02u+2YlAmLlT/v2NXzKxHj0C5ismE
FrYFQSGkmHbPyBCgqWRDJcGq51CcvOD1SKyh8Jp28+gVwHteSv5onAlMRpcSUFz0k9pkWRLHlBnM
1GBsz2Kv8MzPRkpfq54b2ZiRNZ51uO4UpZ5ov0H6Re0rpIrap610TgHK4DrCxOD+VpPOYN6klo27
O/Wt+06iMdmXdKTSB1cu9pRii0hLuDyYrfdXFl/f7AUbrIXl9veSV9sm+egGz/fmWJSPwu4Jn3bH
I3oB4dlo1YvnDE/9kUnyb5JACfc7HDH04/oX10RbnnKtOsg9vDRZ2niP80TnC6NYIu6KQ1Q8WTcA
QyPXLknI38PR+M8psCB8JSP2AnHyoTmNDDXyNfAhOeVM7Klvh2IXM6Y3yZV+WZB0PL7j3dx7Xezq
wSpE/qrJ0Qehw7B2S63jARrGwzyMsVywXnIn/YNq6uJs6SC7YBMANCgGcHCJTEDkyklvcVLHqNEG
KRIIJxmNGCDVfpsLZW3WMGArAwV/E1wleRNdlggp3DB8MBW88L6ClR5Za5w6rl1p0GCXyhmZx/yM
wVZjiLnkp836039JrOy4S5y00ZA1/Z/EQh392VGMmeXECVV4NOyUmsXfQO1daL7bP2QeV3XduKgN
y3MntsmTgbrd4DS977woab2f6KWfxAqzIstd7W1UcYs6jZXXSTqU4EfoyUtPwJUxjK9N1i9MT3TH
Pe3pPwZFy/8UBq5Ggc3FhgCJOw2v5oMQFPyyTflf+aT3QqsOZ5k1L9UT7CnWt7556VpDOZRZhJFC
BIqwAp/LaSCIErzouEeB+ggaE6JsI4UcJ6XdrM0wTALjGfZN+zw0Ga+XJR18i0+WJw4Wm8cqY4Qq
pGsILrV4IvQ/EShOav6hf0xn9tFS2TXXYdl0hIhGMzQ1DQB1yQq3sleudQ7BjedCLFfQEERMdS81
MUEgg88NjpilX4ECnyjPLcm45Gx6R2BFmQkFW4mMrCrnszKXreYwpiSu+cr2Ro1hPA9qND4nPnkW
x9/jm1IPLIj1mvme/4yBJzumK+t+ayy47u8TNIuEJtGtqJXrNfNSYI/3K+DCT9ghuF/06TWjpb+M
6U4La/wzoZVGHJOGxBAsCg9iBPA1lJPryKnCR1L6LX8buCBdT4pFoFP395hmnmoRgaxQq1dRlqlY
Vuogg5zVt7+QFMBZFpkFmFoYCl9qpYDXN3bTAC8OR6LZ0c6HJl8yYHkezrmafPpwACwEgZ9sMo+/
57nyt0Jhn9bXQ98S2MpUyNfGejrcy1gfpIZ5AlwEIcHq+zJxPIcyABvgzyqFs8v3dU9QxQa2Sf+j
7lh2207luM2uBW6AKn8zOufT/Psw3ZLOOKXxiikS6rxCSO8lFEceUqito6eGfYu2hbpfEE3AAiQt
mFWz4ZWrkRlAtMwbJQH8jmwigaDKe2PU6M/17wWy+UNJel14atZvR8lOc6lclxN9DhQyZhvs+6+5
e6do4YFm6GgWdEgCbuR14VCm3ZKdS13vY2LwjhDpmRYBFMtszjLCOPtvoxwxLHjpnB0IgaeIVNUK
/Wrw7qAHjC+LzaYH6m8MWK/5GMe7vBiOBWkeEdEZJIA3mFuPRZEDEmfBmwzb9H5F9YXdEZvGW0iu
DC6QhIOQppE1a7OGU6sfgMH92HkGlBxLUK8/krPNEO8LtepmaUHpzFw4d6aQV2UqjbRdJObP1nW+
C6mA5Jcxhby52qLigoScrIrJ4VMHXWTMAhLIbrIFV91+XUANrVYUy16rcTdCmTyDJCWJbYozkKto
L+aZPDFxmJ0Iim7ceskJpN1ZISREq/5h6zLCfzcwMhuIIefXi2rCJ56jZHZNm9QGaX8jdYXiwp0b
HkNWJFtTiCpFNhV/PewyQvlJpLbS4PjVXzkvQwcX0Yw4FDuOXKMQhl0joLn0Tr34DN+OHJhEWnIM
ar11fzhTXZeYGHnFRagIf5yLkZYDQJIrn1MWSoYlp9ANnGGSCbKwVetPKGkRvyc3NSUfCjE0vEa5
ujgWJq/NklRxaFE3aG7+xNo+O+Ct9ECLfm/2NtSyhY5T93aYCFVEKRSjjeVxOe4bWb4BN6V+3XZV
Uh6SH0PmuNkdhYkhbB3dQFPVDaTHM1PwnX+ninuxnrnpgdjC3NMlHlWC7Up4+secEwrWQ96/T+v9
0uvxgvGg66sgky2IVed0iyc2kEUSpQgfWdEya6CjAqQGYJcr8o7zTmTeHs5t70jQhlPG1g3ylUCh
dGxk5PXVqI3mxf04gR7EqlLNq9w/yQynng+2LU6VpnHxj0kAc3yxlieQsIlp/hi59Z8/7lBnwzVP
j2df1yv9MN60PiynMmQbbb0gLv05YqWbzbf1ZyL4yePescCcvvI2T5iAwGzbwaNMh6DYG/RfgjOf
kKrU3ysHPX6aXGUva6WZd95RYlLV75Ro0czM0Q4hB3afPtHJTJm9qi0B2UbJAhv95dR/jz6PTlxm
1Daob1sbzhzImRBwL73Jj4tjbcbzWQuPXrn4qpUJYGU6e8NuoJ4om+vWtbBm1UFOwnlms9TeC3gw
xCegTl69NK/xlQkvZJBZnvPq+V4IeDYMu5e4Xc1bUybPPncRED65MJCWdSx8llqyjsomr9rEK8G9
wdhQDwTXwKx6IBm0mcpwTdC3YHeFj/t0lsAck5epsWO8FO0H/xDe/efwUxWQu/S/HjQzer4lyTDH
mwtr4Zs2Xjz9Z+6VayJ7fzMcwyEdUtiZMvDqtNjW3BbwkbLCKdvlDPPmunIXDTw1ZTXqgOg88oFP
FsLrD5N7KuBzUBoRtTzd1x2I3fAWIvJMFbYqpjbNyIO+9MeCYqCSOky061PScjGy/h9HLbmsxd2I
xAT8jTvoXRnS40/ia7GxDOtRiUEUOhgFA46fU7L19J0pdzRCaTRP1TxTQQ3mAyPYXaGZi6cI+dP6
YCZPJzOpvxlc9Z45KqJTdMyHBP3zTW+nJvN/3vQ6PdpgtXv1jsTUpatwukxHiwhDBPe80oTZq/2R
glNVwwbF4S5lRH1S9PehH8c3xs5oZ13/tL5TgcQjcw+tD8mLhQ72xZdap8T5i7eWeUkmctPQIsfX
eqoGbo3FZNDt47dleERTJ4KviC+TZc7ksetTDBOUsMnRPmxCWDjhXSjihKVl3vslaEf7bR0fSwBT
jl+ZDA6iUxbUyqDmoTqzYVEzOO1svR690/mY/bChKRiMlatCqKuLHhW2DOXJ+1GO09Oh1YHQW6co
f34OaMNsxkydavJJb7IrN3kAbUZZT3w+KpIJMv9tu036k6pEGOLS3SE7aLTQSTN6Dx9qAd3UNlkJ
VvOyfTfJpYFooTy7UWIb6v9Z5q2Zly+zHT6cxA0rc+3wtDAvScZONDmJx9TzX+fP21OE6PqN7Jyh
8irK1yKdpJi6X7SYj+SPr8ttdJPV7Yxt74WqpW352UTa/exYzFD2qt5Ln+JToGKCQqaw3J3bVe3q
782LPkRH5Ic711c4lJuA5gdKwTtpcxWHJBRUgvcPI0BshBVgqUvM6DzTe7wQ1kISN5PH/3msjcXo
K5SzML204v6usmmBi7pxclo7fX+1xmPvCCpND9vGUUDrU4q+sHZ/IK9TwTcQaaAKJhPd+tPMCmC/
dBQj8CZTwy/5zYUP0u3EXl9IyviNBVWCnSb3b59tDBBljYja8B1Q/uHJPyS0JKa5D0Zz89LVnhDr
aMe869LUKy6iMlWA3Fc415fAUW1FqXPZBlS1d358qQfGMKflCmQHUAbxiYysR4gmCRez3LhVS8kH
9uLzoPgHr0+/Zo0vSSLg9StXm01Cc5DaFp1E261HfiNHCoq94n46llf+gq9JbFAmmK2FCuz24vni
yc3e+0k12IubjvPeTspoS9Y9o2WTebS4PBsAMMJpky7Y+FYH8uTWGss4A9tcJToq4+fp9c8SlqKs
GVjTAT+kdqZFMQsj0Y3NAc/9cn8XEUunx9PITmekniZ0Sk8xcKRWC4b5dXoLQUtxvNFn63l5DZXb
rherBhpZJLgd8Dj+3AwIrec2wtd3Y5jUmYwFROVIiM/izRAQDkxeAWkiMlwpMRnFMhHIktdwF4WH
q+nJQam+8tZcWUSkScplgDnwY28KsyUl3RaB8WVpVUNIwGIsDfaHAMzBTFymSEfTvtUOWdB0uGji
SMS4ymv18qUWIPWLyDNdiGEnG7KxaAJ9Ez1AGh4w0oyPpanPyGvYB3ysMPKdd4eeYVbNYPBbitp5
xpSxW5WlTe7F4yQoK0SL74hVV1p9awXpGikEOzzVLVXN7mkm2tqTpvN/RCJz6Uts/kmlBAousUz+
PKFePRRnmq/U49zuFF2Fc67ATNbKdJ6QZQRm22w0O44rt9dqNnuhXdEuPKVqarAx892nmgcd7CGR
ZQff64dEJGRbln/2vUBdyNE9J6mn5R7vfGiqMkAzjXwn6DTyR6Vf3pek3JO2/Zy/ozHwr6GMuiLy
yWNEbG+viNUw4BdYEGa4fPTjexXG8zwEk/79CJ15XgeaNc9jJE3LjO/fEHtEeOnnhQbKIepcrffA
FTm9sNorf7TU11GKJ2x2PpCiePA8J37HfD2u+lEQrQIOvnQgZuvD8ZHwH5xavRUpXpgSZ1uIrIJr
CLT2WJNI/hv1yi63BeB3wekDUH4/mKEnMaswuudeuNOKOYSILlVvuSTJZxhJF18PJTeoJUxJ1ZTt
VjwqijEf485FwyRMB2eD3yUU1h+bjXLXYydFZFt+UE+Wr0WDNA7fU3nPKr8F1KAZE4fNCp7sh+iK
YlsGv4rNE4pKNFJLwiS+Q8JO499hvd+Bx+2Clw9dOserGauI7yWVy/nuH8FBVvz+TiqF44izT1KO
rZQYF0FPg9nlkHskVZTFsuTA1P3qDRzogQbRGi4r/WfEsEnqx9l3NRxM1r3u8LNNHaq0Gdvu9hyG
mMlfG9NIdDZImIAGijiTi5xCEtqIgKFA1cY5Ot5kZCXe8bgkiOEukuF+3NQbw4WhOgphVhFk1rDU
HwrHoMVqpJj12DvcytJG1KNx3IKji1Cb1M+ScEgVO0FHPaMh12NNLg255TS0f8SRI7OvrL7YmzuF
WDWD3fNF5vhyVbrCaL/bY0q6ld6BceRvntiH7kjH2hOutR4Q95snwRO+NJIByZOZPguuOFrHNKIr
OgXgIXR9tcHQxD/qvbTX9p0108sQjCNvkVdOVP4igrYzvptn28oFtDYqGVdXpp+De3/CHX9L/nsG
M9f02LLkyC3l2YntECFfG2A/lPtbSucpigKFfzu36H6HxFM4xzSpvVx/91RXoNf9AEci1ixAlEZH
gCCUBv09zaF5YzdWWxgkul68hBKV5O/81zppY2z9NBO/1RTgw19fKRVRV//ycTG80kLtNLBnjqyB
2GJ1S48L6lkRjZgpnE5bv+6kKN2k2gGuryYe/Kp/E/lsXpiu7Pi+oQ+4zMExwkZRvfY+qcsS6Tvu
qFsA/eDvuPqExd0NLXLzkzaZcb7t0YIWW+fVeikhr8EcWgn/t6Ezb1CJMtKTEBmPpjLV4v2jZjMv
4Zj2swhGIWlIKqoR4Sv619dK4zwWnT0tliRjtwtF4DRnDFvJQSbFqLYsje1fJOJIF9UEWjNVVKKm
BuzEJvXZFhRvoj7RaGgMvgKtzsBKVQ9FOacyCvG1IVYz72eQ9YuxzXfim7rx6aqilCNnhoAq5T94
euz0Aa5jq3ZFg3ATg/3/twmFGTLTPmbaJbC7w//5l8W67L/7Axx/0+U+kSa/0wYsfDIwqAR5D+kC
qrQ1h3zyheLnjiitIaPuM9u1/b2QA6eLym0sZ7Jwv4fogPIc7IHSGtnl7eUqdTmC5Ua3PcC8UMNp
3h8jsItKuwRMewEJDvQUhm1mEfvIc2uhVoj604IKDxbuGTa1XhyeFtNKKUW768j8+qCWPqcJvrD+
0pFQumw8ALltDz+uEhvTugdd7fSt4ccOdUcclmUYK1DrlpP/m/PMjY5jO0AvqOSWg2LKD4R3Y1eX
d30iPZbpgiEzX/YIeG+oondGc7v7+mQEOYSS1lEo06ZhDQRpX/k7gWUShl0S4TW8wBomknQqGC4n
gQwv7DCv0O56esfCe8zq873eNECW28DDdnlECd9w+jiChS/T3KdSmKNK0jux4W8qUMRdJmnAsvLI
IfYz7LI9MW6g1/scQiW9I/P/rvHRM8VZzgDkxO3t02WGUfMa/C+zw31OVg/RAMbfQtvrjyn9kFoD
m0y6qeabe1D5Hn5qHZ4bi2FQHFwX75g05b7jCp4YeOI3ZLI4hqB5YV7zqgwbbcA7eS3R+L8XLRj+
0/7n6YXO+MmqbktiyFAJNvrvoapWeE/JTqvFAEI3Gt1G2Gcs7XoJ52KfY84hEBft5nfgnYipSFrK
xWKntwv+Qmce+YJ6OCQEdB/N93vFUrGWoESjdYbTUYBRixDToogBFMtCLh+ohIGbViqweFFmbGE1
1qtdVjEgAGT1HSvA7RP61dQwwFsJJjnmnppaiqDIQfrV5e9pO+zsTwnipXaq9UzNBSYdiuxNboQN
vx5sNZHehz/fnTnqzZNVIVuIWDe2Ahs7UzE9k9NfULI/ObXUWy+SAs2X2hs66CVJeC2iao9Y3fKJ
H1T/p5mI9bAGZ9ACqnnX2Dd9FPRWoE1wlNYj+z7d+Que42RWny2IXUN6PUthjJjrJCyzlIR2t4ge
ZvNi0WGgu5eyJsZaQTdEtx6WYE5I1XuAqzi1jTQduQnyDllGlBPzf931ljsRFy6eZ8bsCKYhIRE0
JQ14cumJCwavOy3wBjCXAiTOeLEgeWYC68MRq4z4OT1zrozzIYmhwksnhVMUlV5q45FUf7kcWKlT
znJTscpO/TcZwmQ6PXEMp+eLNYwndPkXT99M0SJlVyoc7WKsHLbwsKwvNP0L8H+QFXp4Epel+1jQ
W4UZYgHDiQzmhAdFCVroF3dO7MTo3whFdyHvdbOzCnWg7fZ603vBg4bhUA3jyAaLNc+0F3dvVmvw
loI8zUfLnfk6Ql8JR8ZmiJaQOhlNEMgA2vDgnCXS0pqKCaJYqhtfz6orejJ1d2gd4kkrwQdu/cIk
P+iPda1gOX6SYWDVnGNC2a0fsQvHm4iW6VDNxtIz/T80ICZvhEByv+toql6WgBYfkEFuNeOkFcb6
IbzLT5CC6abL/6fOWuWeOJZJZTzwIHnKl16VgZ6COAVO9lRY0rbkCtaqigkqQiD8jV+cKDozkVAx
McbfhJPLuLlSKDvAkzlEJ0Y6wX3CfQ0ejQghl/4R12/im9aYCOQNPT21hR+IMbqOw1RyM3G0AkP9
Dw3PrIkho1VYKNJaiMXuERya2Q6w8ceWcG8kRSWmp2i3buTRsqx3xnyWADYi5MUb9RSU/GEhfAPF
grqfBn5fg2ZVzMIxAFHkG7N2/+swy9VCujytYiknSZMkgSClKIBpe6wwBSW2OdKzWpB21+cbQpVO
wHf+IVKzC9DQikeYutdXP23MClf1l9i/jhNZeyK639GLWh+GFUGhzQZ44xdjtq3pK4uoQdhpc+5z
QXX47w3UsE+kXYupB1UW9HBn4ZpQ/FDmAHGh/CUGF69vPdpCE7OjXL4FwhBw5VUQRVomtKVdnI4L
BX1GlAtbM3rQ8up4dc93nKV4clsGzjAncPKrtRKcl1WlCrqySzIFU4Moguwa/a5OgHJAa2VvCSOB
Syl9JsNv8NPaVHiDFQ85jzm2OFc1ENEX2J9JNPfz3Q8aEE632sV1LJQlGZlT4PH9Ke/+0GSFaxh7
k3Ddio1gsmCz730ldm3RKeQ7NRK4dLGES/osYZXbMRFDgVsEKjoTSW1kqFVNzqhDrMmTCeiXxnXQ
nHL+WCDAC4SE4wlMndbnNYAHDxOExh3TW93jEYkIxePl1Q9O0e0buCtrzpZws0fpCvkKflUqKuuC
M+VZDNI5/EOVFs8NhpTmIRe5yKPG20BLeW6ohcEszgNfQD9GbiLRgjGl89Xvk4+gK0vNVmACZDPP
y0SdASrqX9bUwcYSaiXqAflUD8Mm6FjZXspSHyvvVO/LVXIx+S5ImjY0ad24v5x+hSJVta4tSKtC
71/fPL/JTlzbUkwBpLL/RIIdVPmKEDGPH1nX3V1mqx/HcC56U/grHB518NdYCe3wBtZQR8iZDO+D
TD7RN0TfNaps7AEp1wxVEy8fzlW+4/lZTisWnWW9uUf2ofD3wdceqn8zTyLqY8YcnYgr0fFTxEJn
xK/TO1gfuf0ZgzIHOi3fy7FjhLNvBXccmWJXXnFAm7gNrGKpjD41fN6u+tDZ3JAvkBGv8mULFrvw
uAqJ6EIMk7HQwHPeICuJX8jwu/SplGhciIv/2j6XfFSes6T64p+eobNtny+zzGnCouk/ECkQVbKC
pdi4yzR4m6r2+ureBtRMirYvw9bSN7/IMk5kquHpsMMyElmqCy9hSIslDmY+6dwtAShYmjMMs0HT
FtZyHoC1aGyUald5ewHQJ4MXOeZplSt0ZJudHpfPygF0ifssC7nh7W2IwFzuyum06493XN2oZxMZ
zKX0doQrWYIdCq87NC/qAAN7Kwlphu4UV4ayxoJR/szjYBfjKdHbBWC8AJbNHmBOikiPouSoXw8d
LwEbcKapWqz2iL8n4oMeLjYD+SoEIZ/MMJyAzAmXospqrFhGFpfh7HN3xCuh94MxkbV6GTwyHReY
HDhdjMV+AZXx+dBmJQcIY5WzrD1jGOWkunOGkeC7+xGjZIDh6lzycdPqXJZ+SIVWmEKw9uIuRvBa
FqBhPM4hcvh26R1jqBSPInCAuDbxkdLNUeEscr5qHxfheVnN6dXSfVWOrfdpIMCjeYhVV4moRwAZ
tQKmbwJ+k83gUwLM0tHpuooHCqJReaJcCV+QK1S25QSjoii1Lh5fLEazLUDdRp7cUes2DpAX22Tf
cMyuEaVzMrl9mBjhHlFQVW3WZqfWwtIjKEhvrsbvZBWEUYU15oTsiYpkNnfEN3BNvo9lPV1cVlSm
Fq+iTjB8X/DvLIFJkYPQX1R7VPdX64LS4M11VJhUU2w+KQTrNPSXaszQj2oeY91mfotp6Llq/xTl
hP7PNEu464Oht5v202BeahgEqP6BzfoASNuStcfHqlcYODofxUV2rcdixHM3nR3XM5Iiq8JmyVFp
hbBWavg/msVu3y3iS46x02HEiRRszJ/RLO8La9f6nk5GMyjTpJE3Xt+d2/uXtvzbXu7UfKWzpwk5
mLknte/UWkZ6qAXPuq1SYsk8CQAEdD9JQ/+Hr/uX+KCUuLKOz7kFfdqFo5pdhWS25MtOKOOJAGZ8
tr6kTFjcxo3MMBbNGh2HS1valqMkCf19aGEMQ6qyZctGzF93ZWbqfALX/Gk3VAFaAaWs8WrCiK+B
b9YXp42ID6cQg26xnuug6z0JY/hFVxAnu9sBy3kV1KP9AQB2M0N3yhmLZtE9/pgWaPudnnKMq/Wq
5vz6AtY8qN5qshR0whZ8ngLbCzpP0qhYQ+BpVvxx9pqqnNfBDONDSvj8jV8ZnW2xsHItaiHkSAoA
dTsRgOovTirZJD/A3x77/cGLKuudzVbO23f8qHsBewmjKrZQW04zx/0MdEvo84TKSLBkphKs5/QM
gMJcSI4CsyNwUPVNkPLlNOhbqT+o+gmh8ZzqXBFtZYG6JqcXF23sqeJZgXzAEdwzvWbZhi9XxU2Z
IK0447L+KSv5ZOrlosB6fBz/I25qgfnUdxpWuM1iVw6kqfNkX+P4us94/aegpeui9F0cQay+pG20
nCJ9H3RZ1aFCFhiHmLDR3LzL8s/0nwcy1RoZLhxBrCIel94bY6dFvItWUOe7eplYeUoedsOGk5sd
Qhhk0X8z7HAWmqNVgnrm8NBL1TFDu+i2pgZGMVwwmDrzcPQC7vRp4lmNlReDQPpncl5gH10rkUcA
LPnabbrClHZ6N12HOsF1Asn9H1H6DEh00/SwpXv5G0PlUC3f6jt/Wvcc+BfxIXVmIt0eHJd0ac0h
tMiC2n/wz2v6vjV/bVdIrCcr+w41mHEaINeQHAsK0JRPvVb9BbCermjQ321KR9ssF/1HgLcEOQUR
JHA8vYlT7PQhNjChAx3Z8NJ2omWty/fjOSnMyKdG7qeC2MbGDgrBmITA9MbiyNU71WGApn+QJ9tO
25pdEKOG7hO0SlCSCns7j2YS4fBERGuBTp0oH4JrokCy0Rx8edvjvVfzhyAUJ21Euxvf967CqOji
9zlYKAz0zk+L2IL8f6RajWoTtFyXf99c9QjmpwkeJ0NtBxCeMOHxhFzu1NYLst5uk591m6ZxNLM+
sUqoRE7LF3Axtykr/XSUiDE3MtZaNcD+xwoxJlZljAon4BsEBZaooMdXniMYNiGoVHSuKPSnOIDq
cBkfQHUCoJBMx4yLZviX4pvspnaVrQo3Tu8nr9e9ea8VoJNcU9Yod3Yoxe0Cr/dLdcK4eFDIgDHp
kchlTpjRApbRXIMBd92zLsa6ca6dfCRTLKralevlp8pjHBWQdEPqbN+c//RuDKSfVEVNDxKVVv9S
0SP55bl/HQySTMew1FBJxWQywVQ77YOi7+G2VV4Y1i1/CtCNh44l2rR1tbgpxQPvmJhllDTDCcjO
xz1FpttFq+wAJRGvzO+8VnLoNZoaCQ76vLt1L/iWoux94rjGQb8clAZbNHsQ5b2AZJnMReeQdKsT
5Pm/TY9lEgBl4JMSuAl+07iKJIQij7qVuI2plKiiJI/bxEGeRYKeW1w1UMSL6F56RGwOlj6yxAo6
is8/ypg6tXp3uraImpwdljD+03v/isHWy3gFJAf0rIo6ln+Rvm4MtC/pcSuXfDREhD8PVucCjHxW
sA8iVZ6+x6e5+tTdcmGLfpbn+5ScVbUgumMljzYWKjS6TvhMU1wToD3IAmgMMkV/yYUjsOnD4W7v
c98bbx8oJqinjbh51rVQxXSd2/CQx3lA5s5BvHykKyZoy1QFnxDoxZgjf14CREAfpz9EMEsO9Jyc
SznF47Av4QNg4hn1YrhHfpLfGuO03VNOosORrldYPY1XkIyvMIIvis6+UTBMRhB5AGgzadgFF7ob
7P3p06QtyK//NBgqKuNglxoq+/3MNd35l5s668uxlQ0e+w6+IX/fbWD0IBVEKM5SSVnNjVIJNCL6
bnverjqrHa1iN9IDXyaDS4DZ2PNSSofTicHYbQT9Sd5RLQWKgK6vpwKkKaD75X0+w/N1WZzJes2h
BlKzxxyCOxY30A/njik34Tw6KfLHXQ/FpZaRYlhWsGUm9KIRIHXtH6RwU9pPaZDg3WLrawr7GNtV
HAjTGXo+rTQwvEc59loizFUf9lUqgIfn2Bzxxb8xYpWiLzpR7z73AzkzddOf1FRwGAZm+bTTn+GE
yjfdjwPurHGD5yH1TooU/PiPdb+71RB+jSOwVBmxrmtFpn+PQCgLgZPAyMbhSq+jh64FiBH5u0Yc
h4AY7dWrcoqNmam8JjJhQ3bOngka+po/fqVP743gxm7BK5+CasiZnJNfMtcNj6N5q/gFUeJYLdWV
o5aqJj7Ce+Mkrm8V1sigVeDG8PdKmSUk9uaw6O7snZGSdItILw6EteX1J+gsN63Bt2ZpHnf5j1mo
OhKMwcIGvBw19XEOPz5sEsKDMJKzQMdSvbcREM4uziOIB9QBFcLq/VJ8KbeA+cVBxFqp1UQ6JLV+
zHiMy1vfHKeGp8noUd26DozamoCpUUKo8nqF1bpQ6/IGNKV//CjaL/9dEvmV9VltwmvTg88JEuSI
SF3PGmEzfXRbodw3ykPOwdx5VE/AXX8X+G3j5DPbnL6+KJUcT+Iv6FWbU4dLJaiH4Mx+sOrvX+Kq
QouDXYKSh9lPsCcRLWWgFVuBRObRjd8Bp+CkSv6FKPwje2gMRiBe39+etazsqRJFLXs9wcsHkz5A
W/azfYlVADZdIfNP7m70zuaziH0IK18X+uL/i5xms+3IG3aXncScvRX+KjkslHTfzPFhhSynoF3F
iIP/vcCkm2QfEaDoznYe1svttDMEH2/U5hwj/jIdClr5r7VI//8LHTm4wjf+6W/QfB3KLEV85C7j
GB0FIUkzD9gVsNfQ0EDi0DjABkfWgc2jbnDHZ2Tarfvk/q3v2tGlvIQpIe5gWbE8jiA0o8565ieJ
++SZPTrAMhw51IriaPYpebWZzLy2Iu+URVLzrD5ENOPmKwqUoT97OwVAJaKbdrhVI61qnD5gexgV
+2NcH6/E2qA8N1syaCiCIuNAAaiZtg1rUyo+tTdCEYu2bs+/pduW1WIXl35cTs36draXl2zsk4MN
hZJWv/nM95lmaH8j+MCcnXjnQBPmnvJxG6kmTDNVEajidd0GZSk5fr/NaJoXpYpwDd1NEZ4WKDmI
ylh9+2Fx1US8jF0ogiSCwvGP+2sQYz41ktt9vhthZo3bPNC/F6PMWRjNOyHVEkpVs9hEYeKgMIfG
aTpvMcHnMmOUUbmVky1/jCBNu1A8TxPimjUeDlnVQezOgismqn6miP8zcayiRN5PQ4B4XwqzAStn
qBL3H9m3kj/dX9aM/oSpSBT6iQUFMt0TDHv/7BcaucGdlws4qtszantt0qaRCn2SfcfrzdHzMLgd
+uB3EhCGQYP7kiJnzTu9fXR9Z95ytoPQhfGJdKmmIUpYnQl2ysy9pYCRmtsYf8NsMY2BWaa2fLat
tEBCq+EPgaIhn4TlqO4kwmgSeAdGt5JbHysJFLr0BF3YiesR6vco/jFHyAKRXVn+OklGTRZln+Jj
pdktqGLuhNeXBfDgrksLwscnMPK2meE8DOgQy+Ie927ViH5/FbAdHMDPHVwxpoqIVSoPTx7rzSGX
xMy80vUVhAHaWt+sldaAaDTCJQIF0lBCGpxfF7iaEhT76boNU3EU8Lu/K3qa5yVyKSxLOwrapFXj
lmMPPX4JQaJ8zUvDvytq2cVyCeMemhLqvYntvdB+ajWlQUxyfjzy5+hULDWMpr1UNSGUcLpoZklj
rcqoeMKMlu02adefJP7hHzFzC9A7Z30WjRfrwR+/A5B/rMkQ98WqzUXsDj/jobvpGk2g6FqFqxhn
UC5F0vwPG07/CcfAhZtgCTnNeXcsZKIR+KfLIg5uu3MUcQYHK895KoIaevYjIn+4BYt1y+9HITYw
axAjEtyDzu58ACN84CQPlR00RXwWEssA6nTOn5/Xplw4ibuMT3mYJZoF0tpoaVl6c7xSk7ICqCnu
T35lah7gg5O3W+mrH54TXiJS8CkNJf3I15P/s2KijgpeZo3g/PUjdVMw6Vkes4IZnp/8LUMcKnTO
Yd+dizgFZsy6kNNg054AdzrlpuHvF94Ss+58B3ulM/ekjFJbgVcjtgVD5kjWyyMiNm61pGNI49OI
6May9aFiIUU4xObgBLnOllBbwr190UIatGgBi3EsPVITEPURU0sk1O4Etlzbz2IssG6BUtuhhO2c
C/ECk7uZRaiCFRpHbB3kINcCgi/Bpv8bVmJP+V1SkD3sIu5YsIilwrWhi9D/WjTFG9NiKHsZzUqE
quPyHAgTyWA4jiRQ+X0xQOgDgQRlsu8B4k2aqbUFtQF/m80SAZkH2HpR9oQtNWu50x/eR4plzcev
Evk76Vbab4yp1x/ssCjDD2aqbrbi/za8XYQkhrV7PER045Wq5UyztqqSDaKJjSTBbuqSp/sdYSnq
nu5iECSXV3N4eMl/taopKsz1BTRkRwid6k0aLQip5CVGq8FVx03JsnKBbZErl5afc8F+/VUqqpfn
ouBEWnLGmqQdQWZd2Vx9aZB8Okqu2e9hu2zRLN8xZTL40vE2sN0WgAE2cl/c0mz9ZBVIVLQ4ph52
Wp+UA/SuzOL4stT9+RUXvw48qWVl8r/yF6ktwgk0/ZZVlr/mDGCfjJJZPTwV+Q3wsYmRkSG/WS4P
xeteJMZ4QDE+b7kbUKMtBGJJrFq2CjxEqC2fpzYcSexv2HmfUK619MQWtuSYFyCXvOmDPnqidxAL
W+NbIxBXzQtFMx2fHldRvrosSbccNDasEeFdo+QcodHAEopykLqalFMolw46BKQV7XTAX3fxPqp5
2v/qa4nrnyBjFt+9/5qBycatAxAD0kUF25V+nZiA4iJzS8DQAK7xdeLxQiFH03UnSsOGCzvmhi3A
EeKBfFaqQ0As5Ck6YyEVxFZo2qofg15CD/AS2snTyHhRcsO1YBKon7Lf9vrMEZf56jctcGZy3d/z
nH9OC2HAau2HjNfSsVj9VVi/2ISY1B/9Ure7ianyJ3Be4KWvCpIiJgClI4np21jQaw+ypXH7bhxZ
mj4+pvoySTuBOhYs+es0Rcy8BxCczykqluc3I5qPpHg8dcjfq5VvtO5s0zsieJnPYgWWxPprqig2
AQrGO059wiJenJgDJkrZtx8JENVIk9gEF7wXOrt9kPvX8jrsqtP9xX0LtQ+rvOr3PhJap6DO5/dC
YdYvLYlFeQtm3Ml7lQsKIg1a8YdiT+UEV1Yzm2PILK6D/IjTgU5VPKXORfHcD8+V7m3xw6QEEyZX
Qd9re+VTOsjSMr+oxw/0F1oxqo0uur2SWFVTOK+JhlA0FQgWGfMCSApYe6kMdt5I6FcxcjpyJwIA
xo0mJG+vx0q5DIwk6SyQS9HGhMZZ2xCPZgu8yDenwIoEXb8JYAaFtFSFBy0CvoXRGzexgEL+kees
1VbbFvFGIsuQ1mP5h6aUBj1nRLwMc48ADVahuGxbegf3EoOqh8PEHYpTJrII8fYzOvFBfiDlxFvh
dX5u7Spcy3k2rm5Cd8cjLjUFjPjHw89SlKWBOH2UAQ4t1+fsS37Prq0TdkVFPTz+h2XkdJGnhjGM
w8RSD7+NkPDsmgTcONkRB93ksn5AJ68HufUFR2HaaSj7rG9HiZKJypcjuA9SNzXbgFML89QiLl1d
9kXUgPQ6FWzuhKhIxH+mQMkLJw5iFcHxK7aaskxuGB8qemG99LHSzgfrMskcWhwJ+Ba4PR7OlH1a
cu6XIvdOaY38Gjsz5ke4AEbyFERsLZjYNMKk5bhpaxFGXvQAzhKRJQ0EEIKjR6KDTZmqt+Wasjy0
cTe2UK/oqJuyLXnwklJS2NPnjZDRurxKVKCO5tdtfB/R1cSixW87HcD8r8MaPewmQc1ooUVY52cT
V8SerQ7r+mWeb+UtVqgNtoWO/YqEO3IyRc5LS6WueCz2uJadrSUY0WqC2Ij9nfRKQDsCRLihLrPH
gqAX+9VmalfrazPUph2h0aLHifHHqCcbH5BhcLEYvjD19E/49282ePI9HfxiOwjeS1kd3wzDofus
6Ka8eDnIvup2o3Bjg7DoJ1sjFBfig1dNae0ZFkYCI6h5lf/JzrEo09Km3zRA6b/h0xbDJOw6xNuA
CUVPbZ4bLzZiMAEB2PcchMfjG1VOC0pCuLkmMKoKGdh4ayLpdnopy4BQlp4v9EcqyqNsgJtWyvMx
UDS6i481uh4/TEidllKHqE59lkRuIUoEawvsezHaCaq8OPJRpvJ8qICdMyx+TGkV4IhJE51Q9gGp
MAXTNX8FWO18208PQ0oHEgh/MCfxsXijUTQvXNhjWWoRTicjCBQugqS6lrw5RJWcAEevNRg8vYbR
A6MEK9sUHqzolhXKdTrqzCmPj50hP+9jIbNB0jiws9hrOLmX68HW1ypfTYk/6E+AoRvKU61KbWbX
l8mpdBgRqhButYnBe+2/XDiWjtduNqMPZePWRRFUJkpF5Q+YUoNVm8ASayNQqmknFHn83qPZgxlz
kqwfuBud41GNY0BvweEw+GWpwUy9nsu3BRmBQE3eGReFDp0xAkGC/mdsewBskfubm7O6etnokf0q
6jqmCb8e66+cjXqHAOIsIDlko0MC9Kn3j58ocFI+d1/mRXYHsepAVX/PPmSX8jqs48JGk7fxRFLk
3M2vvZfTs4NIR/y/4amx+49mt26Iwt6NzNKLnNELugcYW65uPlFRc1kzJ13lLRTtrhBjL91ksNbz
E68m7GAH6X4VZC9+KUy3ayojKZ7CS+HdT/LGYwnylbnOFzI6V9tFI4z2sVhpF3sJh1J1UxoW0tRo
lLF4YFeZtuOQ/pXb2adh1Q6LTJhfWvh7wFtKxSqkYwlR4BwAOAAAn2ljUnHaWcPw4VwgIMLEB0m5
tkZ3F/gYPFulPwk3MveffaEv4ToriCPUXnQstOsRxxLl2ceIIdXpWi1DDL4i08FRnWPFAtljftJ2
XMYYsjR/gdB2q5wT12mGOu4lHHEpQCFceV1n/H/ZPYJUy3ZKR7EHY+6vikZl9Qjc3VtU/3tVMuIs
QS8djcWY2tAqzLZeerRQ05pgs4ZuOBWxoJddgyNxgHFhns6bbkjARp5ypJ02jbEr26RFiRoshLUt
MIpxhSV2KAt4vcs/0j5U0h0waFknm6KdjdU7B8netDsrsi3ySVBSgpxbqpP64yJRhX1tHJ797dtz
nqPLBwgdtGTyR+ke2LRJAuq2vZr+QqrsC7LCxdl3hadL2oUO/ZtMe5W0ms5JvXG8LLekuOrtkebQ
1jhzXeHRfHUJxNzp+wd6FfdsWcqQqFyP/Ks9VJmtu+EuNHfWBNTbmThI19iEPyAoAyk/nRqbpHY2
R7Ns83qZ4vMMBA3xF2a6f7uVUvu+Q/G2EPgir+iCp54dVfdgTHWrKXMDKbRNtXFrL5snDD1N2Y+k
Tfz3G1X2SaunwZZJnIL7VKfZeteoCFVFgAEYkR3lOI6I8URGJ26TIq2PghPGXT84sCn2Bs8Czn63
j7mIYNA+kTpbHQmybRDX2FnN662+3or1sIMxD0J1QPgC41Vl8oJeMKoQkFoevj88CsE45WD3IlCM
GSCpJKGB8E68tDp6skYojhBLwRuvw2SgWy8CjYR8Attuo3xqlElXWxlcK12Hr8EA3CuyynGQrr8K
T0n0OyvtyZcL6mMoog/ES7fCxfRi6iolMEXpLqaHDr7o5P5QfKO9PoaS8HKvRmy2DYF2h0rsY6zb
0PhtFayAZUl0y2/AhysQdXPCM5aOh0yRa+QCKStpMcVZuEJUB0bu0mWNMtYRGF3zM9dd6iWAbCWP
3F40ECXsm81EbRx4Edix5S1sGPRVIC8yU2D480/X7oZm0PE4inebZKNMoTl/ueU3xOAi+UAKywqJ
y9ltYHAm8WDA/CtfZ2NJs96igff68AF9qkIilp7mz3z3NIQxJPmgH5XTi4s6tYsbe5qkrrmdqe8w
8oZosqS4iX+pThB1bTLgZAzdCw5kv2E0FfTf+pWpO0r1ek59fahN2/kAyY7pgFHEMFfdrQQqv68s
DmIVpYzU4lJITMP6Qde92BNeTWHDfsNSegz3ky0gwOsFZMLwk0I2f+fhlfRh/WlD5AAnSjSca+y5
2KNlHhLFauc9aZd7tppnh6vvouirCv68pXDjsPlzi0fYWxNs6B5gwVlfEAAH0Z4HGU1F34C4rSEG
CbZ1ZTmFpv87buFYdeTt1YW933nLeVSXtOJLI609RklGZlMQknJp33LPcISLUG47BNcs3KvyvFfA
YYrKVL/jU6vs7cYpAY75N/g/9kjFGbKNxor6pbTNQ8TWCdQGxtOTPN15MECS8y0aXRFI9+GQzecS
2qe2eHXV9/WVOcPT5NfNJiK6Fmhk9od6c96DiZWqUEK6dpkDQBjJsuybHwsdZxUvQ9nx9iq1t49t
mGyrWpu64Y7IFllNaLyLV/NeSrNMqbMKkeVv//ZZkgDuuf3/NPje+G8TNnaPFxso9TnSp1kMDzV1
qS3SBZGgS2iwg0PB0gW6Ljd6fGA2R8xeunE0zcg62bTsP1wtCIXWpSY4R3AFKlWECwqbcxrRxF9d
VxXHVhci2sFvhpIDfYk+mu/pa0GzXJEaMjuE4KIM7QxpBwrwPk3qsNJytGZgu/aJ8Rf9ANpT7RZD
D5RdHFffpfJSL43m+wqgoGFX0gv3VZE8KUlapSrA8Gm4wA5nK5esPnsvs+/s33uCyJa3C0WlHWjR
Vyk2ecu6QE+X6KuA/Km5A5PHXcGZ7/IpTQkhCH2rusJ3JOMZ8tIxXQ04+LeujjQhq9JZ0jGdwgoc
CeHnaAr3o6diKCUJ4ao3HjFREMAwBxm+Xdb8hVpad+B8fgaP84GcI3AKwv09rxFZ4Qdb+x39YKQ2
f+jUBTbSQYW2ltCoBCm13VF05aV0ZKgtx+ViSPdJxGUk0d96w+VQnatEQFai+RsO5G35eejX9ykP
B5M0VDziyQGeE99V9uOIHhVBvY5SLu9Ld/74zDbfpU6HVq4CjSw22DxnTOgbh8dAbio/hmQMES9d
bnavArJds1TksacF8y4oE2M+qVjtYx/5yVY1yUgdxSS7dK4Y0bXhe5CxZJTvJd1K1HD619zCarW8
c1Fjw3sg+m/i2hbXKvepADt4JiVV0qgZz6lNc8ZGVWdqZKXxZY8ibU8+iSOaTlVMFEW78XduqozA
uYGOq7d5gla44pToENgY2LggwnQHoOnPq/voQVt8YffLmlj059ZOVUtySgZejeu18EizSBISLCKO
Kh+sZuh5UeCew7w06xPDLZTyiQQ+riog+PKfoEfT2fM2bC4Pnnxv/g4MaJy2UnVnZc96kRwTT6Gv
Dcw3XrzUx6glJk156Ef+DyBggbIt3s/3X6IJYb/1XErgWI2o1rXiDer2oKzl9WbO40bQNOVyRfjx
B0doHkOE0g6pRVcfIP1PSg1WGW/vWToUy1MEnUf5qaFIPHgmsWdV7I3k9rSYIw7d8c20g/aLgQPf
jPwZaNUSXra2zluKEkLcudm4vBcgpXKBBgOHQGUekn8MLe/Fjbiuj3Kpg2n7DwjL6ZVi/BgIF/qL
Qi8ojwiBwXtM1K9otrNRdEhpJQbyrOQWCrMNXjSo7p6hAkU5rG1K0tNvVNw4nJK4I19kiytqeoQ+
nSah5xX7MnrbyCaeHOIkqYMA9ddFwqyg3+C6LjvQlTKmJQygvyk+FsITTJ4YRbxxos527WhU7OIH
dixGr29l+3p9SKoOImNY/VBwFmcxF7Od5GJGS77ynT5e+xaVFdLONZNmdHe6WB9rEXNz1Y6P0zAT
4imtzbehLxFpc2GzraaFdVKltNMIk8FCj1Yog6htX5hM2xtr666aLapkc/ug6J4KYXt/0H2OKMsk
ldIqW8rUXCQz4YVpRqIU8818TI8KXPZ0AMh5mFJzgTeIaQx9euAFF211X/V2wJNkw/Jzgd9jEgoZ
T0nUQ+pS78Iu6nTDF1f1glsP3wwwCsLEbJwa0sZ1ykUns/Gt0x4WtCL8pjgKWFc/kIdOj5o2VsQj
OnlTSDWZWQ/C5oN1lp+Y7iEs5tR0+gQwsFey8+9obPEVVzc/sf1T3WbdZfu9r+NsVuc41l+xRAAd
JQzzhIF6z6/VPYdzUcOz9rV4XqD03UcMtn4AEtD5suoo188IEj5bNyqC/cImaZpZ1NaHEKO3X+Vf
bGYf/k9yvLLOWXiR6GE7/ppAlWWu1ENluko0+S2E6dZO8E6tre+7+H7JpEUo/gYX4S8q5nL1wntO
FYh2L+mPrtL+3mKffgPiFjvJkhmqDRBHe/Tz95bVQFlsLFntcrn1NocUvY1bPo8ZtMWKzMt4RFik
jg/w03oasXDSY3ty85ymyl4tu2L4O/SIWMe/LpCScof7ZRm3/WNayAmb5VB1ROKFKzb7X/sipo24
wdccbCj0jglIUaM4xqir3bvnpkMpbaih2KIWN9cHHBir3+OiI4iK2txHCWmh5WDxtZL7IGYueVjr
Wsholt1Xt+tZ9b9/+sQFsBeWSFIntqI9P2P9IBD+2vHK/JyPrvrxM5Cgdq9RisfOAPX0X1zzVN/C
c/JHn/I+y6+CXNivVzarqgQwFedwC+yN5d5xJDGBh2ixVP5gIL8/GL19ATom2/aYeFaIeXqLmHFJ
pdPgXjYbNawLL5Hxp3HvcI7iMF8u5jUMGqvfrUSp0yblwNk/KBRDilrg81grS0v5diINHxq9FnPZ
yJSuVnEa8F0lY5cUKC1TYfDqmadizwfxuu1EeRK7w43B0BSLqtiXqi2Sx0utDxAyn6Ow3aU+BGfR
p7/5wIF193HSus2aWdfJTkp7ieykfGhcd1YQ84UUnOV2MNusZM/u7VMacDqFR67mx9USGaKv9aql
QQUI6oOcAmGQXDQfu0mgrqzagOfrR/vGW2QmWmyzl0l17yWpOfA3gZgRyG7Xj8NSjhf653iIuxAX
1ABgr1diRziKP59WzOJ6/G6JyCXPIP/xe++eVqVlP9tbnmuymrWJn0YnGUOR4ynB6XCi41mBM9uU
Eb1M9duVGfLRc1/2xIfoqJhee/VmEoZQWWKAISFb4NpPdJM2z1LZbgl0XeN3oRDuLonallP3bJoY
hnGJIjcigEVboZfhDtrJAPqxpkNvuuAM+WyJDfFx10wSNOpg9zEJuLnrYYCVPTTI3XOFUjtTyzs4
sjP5xINFBI0/amMP1ZptRMnKpzqMVxVNGqxGlKywa+xOO5RrS69YQS4EOH34PM/BNEin83k1yHp1
yEpxS2Ur6gDNEQWq7SeAAOLUc0vMvHyVtLwRhlxqnsKgBRpuRLhfTjWsMrdHtxfdvh0h7ncHSvPO
sbvi64Cla99CDYN+4ymeAwUBJnfPlysT708s5ItB3j4L6f87sd9RVDrF7F/wUDO/ErYQ9d/UWN75
Bd7o16eE2bFLNWSQeMLOv3VoecPXor83PwkVdZNfE7mVRdJwEVWCbW4OvtS+rPnmgHraQxr6+AVE
dPv4fIr6eS5N6RuDkqzXP7WPQnpCQHQZM8jVrHX74X+1+ImmsrCswHG/BMlDLuRcjkt+SaIvw/JO
/9nQs5SkAaUsjUk5+X9gSYYZgJS5uSBTFJd+3L3eKAIwsq4I9RMZj6RN2zPIITYpiU6qLoWeVT5P
CMtSCve/53+3sLeVpmvNq71H6iwtV/uYgfTpZOzQDFjeTHTBy88oMTl05+HCrF0hyG6z4lu9E5Ss
k57PY1fk5vHD5n4uUvcNiI0CItVsm68XNcG4rvLJXg6DIADnwG52WStAFFxi2lY23wORPwUCKDg7
lgKqkzo94nPOJKrO8JJuSJp7hIcXb3xURIaTHL1cMcx6qA2trSE0mNTBy6Sg7+BjshWMM/t0SkGO
LIj+y5swOm6MDZX7IofrC9s9vlwCy9CH4PeaKA9CjBX4Q4XGc6uFf6kirJ3xZ5nYNCLc6pKZX4d7
qohC/Y/RKtpriAAjYSsH+GKj8IZxQ2OfK74SZt0IjS20ezWsIDOJgA6ErEqTJJHZ+ePcu80zGKQ4
7ktliT4RmR9fT86pOvnMX0LapjNsdKGU5slVXvMz5XvICKuE+Z/ujlwth+tZPUcxupdY6Vpz6IoM
EmmfmEBx3s14zzaXo8LIbRLV0n1mNr8HazK5R0m6mPYjlUp0e2559VvTPoGT4FWmqkg1Mab0j38G
1ote7a+w8eWs0/9R3NtIWZFzhXgpSOTfgiZQ8YoZS8Cp757yBhILyNV/UY+1A4omgl2alrBlFEsV
w1CC0TiKq2U/oAkfOUk4idOqVkV4YpVc11hNHpVHgS/vGMtGhlPG63CTnB5n5ORQ6Lx6t+auJ8Mu
qGC4uylZ/lVQlCadRTaLIVbdUM0Lbf213cQXTAbZZ66oo4oGTBn/q4KiAT2Fja1UkXvm3udnWY+O
9+fBXH5IocLHsk34CQ4x1F/V7mNgjK1JiUu4waiA9aJPTuzFRW39nuX3KKr4td3J0baWVrKktOIZ
iCCvjziEciU/51i5UZRCGvjDuhIkrgFBFB4rt3QBrj7iw1uvh6P36+VNF2+apccSJE6eyNJB4alj
hZS5czlEynaLmQgPSt7BhaAXQ5zt1ZMsPqwn5Gxx+arEfmMnu2gyScRAXi95v6rH2x6IF6LAOJJn
MXTo9D/DP2vVWro9wisGA+5ZHQFdeDAC/A0zzjYwpdxJiJH6QrLpPzq8WhvPY8YOd9cJUtPqdOrJ
R5AoLTc26XEj08eW/p/HFGRKfQyHHZZy4yq7/Q6aTheccGXotiDiHWmUN3GlyiqcCSmnmLdL4KA4
q+vUz8YQqtGHoEaOmQtsbjS7jG9aPfe2bc5La7pFRSl0j6us0CccseY2QPaxYWzPHNtEtEsahQDI
eiFRFM72hfn73XZWT7nkjvzGQZbYExVUgEInoF32CIqezCUq3H6UK+h/vA0nI3BC1CtJbGQoH3bp
VlYbi4MQdk9mXGIw5JgC475w+Te+caGbAXTlNLFISMNRhv8e+xv1hTKLm8R86dv/VTPidLCyEywq
EHrEXfzWYnfLpNwzsSXFXzxWiTF9YI3CJyKo5Q/BWaF8694f44opD6PCQTAIhBYfJCSJaQAiae9k
q2PYCTJXyVDysk/jIfj3Ufib/6OnynRkJhfsZH9RJqyjMAAbi9HDbmbAPu596HgOslQHYNVypCZK
fLh/B8FQCoDVGDJgUPoauJo0pmDpoAwsiI9/bYNiHPo+FLxdDNxLHwWq45kDN0XFGCXtFXerR7yU
b//jalC96MQwUhgFNI43wz8idWKNGxHGy81ERhamItFPcqjQ5XzwKl55TAtYz160YQoQny/xznew
1TI88RXFtSs2qxYzyb8f6zp6lT7+/s+QQrZ0s24D6oheDQpKtkKqtmAwsBWJbtZITsiVr96VXUu4
Fo9fnM9e3+FqFaIcJ4eZrzE/P/PCc1GWWOS8NmM07qGhQcc6zGf5/IsEPaZHFRCE7mf8mHjLWexH
wAtYu72kZzZ6c0v9uX7/tdrJqV1dJ0dSqdArxiVkhbEYxF0fZX3SbZN01uUIRxbSmQr4ZPnwktK5
it7d4dYWIrwesdU653XkaNUbFME5WyPPoGFSTXcq+0YhrAVjTyyRmgb85/KHFjlA6JAga+pQI+Y3
NI+TOvFl+4AoBnzMc+w2PDXN9PhGfja7gIlJTNmIDskTqEpXLYPa3ZABp9yrPCc+rXe2C7oxXXzb
XbIgGy9ehK3E9cO4qqSeBqkAYxPO46+KVp/FcjAJX8AP8zep9uFxGo+zPK4YYE8DTxsq7tFlboJP
7csHf/lF+Zkqj02zOtqDIZfNmzx2ckkllLBSVFWgzFVw+dGvcUQlTUF4d3cfRcdUosNNs3/J4c1u
ecBXIGJNPoTKfxeF6qHc94FSjAI949YIbRBg6QuP1uKhCFRoVC1z3SSxcsIAYjZbXNot0AiCl7zR
mSRjpYUUCVefnWncU90KJ/aTYQn8n02wqMadyS3QPdHur9nFAXqgnpl1Z7JjZAV/q/UHaTLOiKTK
ceV9OmdaZP5vfZP+ccswWA5xhED1VtBKoLLdh1sHYbGYMzx3AyDNIpmZ+RnB6Bcz69ciOY9pLH1v
Y8PfRe4gNJy7nB9lARY2G2ih9ozaas5h6ITD6GyMeaysW9eFXHMRYIBP1a6z1kviBO2marrTl4FL
ibEozCvymzaYFLAWAnqWWRXYboyN/qYi89EJqc1jctsrxlTig71ozattoQoCPCR5WJRdnK8tpa02
op3/iugVyIDhHqGP+qc7rZAPHZRHHEB760Mcn5n6shrX8olYypDJUXOeoQKyWjLkjMD1MHllwUZ4
7C0saXsZUo5cS2KG2alyba2Qh5rtMSDgdv7YQplbi6beY3mzLwIj9P/idBIaSGNZ9I70JU5KHjfj
1IC6g7awB4HXxTENHaXK8FaFY5IXWJqWa5fQBhpT3fGUGZphxtf/kT3j6bYHZYfLM1rBYm2/216m
ZcW2YzvFqz+J1YV4Yrn2aCH7k+mILaW6WM6C31Ief+8TvBsEJzEr9j+o65ym1Ga8pMuewl+P4vS5
jx8RMkItm5Cu/bzU/c7FabpnWwoZ3BQUG2RPRV+tQw9UUDQv9uQSRQvXv17hG0ndfl2Q8b2sgaMA
c67Vy8Uae3cbNbNz3q4t0V9DcO04QMujhTS7FVfNACBb/UMh5NOrKIu+wXtaa80q3guXkbpl3xf+
PAHgJ9IVpNN5KBwtw02fm6KU6HeLCesJEvO0XQTbLVlNP8FtcPqyYVY51O//vA1o2uMlGrGIqpW6
W1PNvPSl0z2zooOf2nYqHgrh8RvoZHxpF8Hai76bSUvhfSVsVymLR5+j/ls8D/3FO0bylHwrFOor
ZW8sz1RkNqNs+AZEmWnYMZDAYe1opB9p7aKdmXvRnvb+jS8Bd0fAT6rEBscJ4lTKLaec8HJC/xIr
HJ2/OmdCOdYxM2NL/qdsCivlE7TPxwiJZvGGzh8ChCSwpaqHytwk4VjPPT9sERqavzRecCHJYJKO
LXEo4Lmlo0LfTkRdbdiaHVpblsSXdbiudtzvis7T727xDXCh43GSVWigiK+zN3DmaPvwez6R4iPs
cNV0RQJCFZMwlbNNtHVkqFZBgeEs8NX5GUAWH5TV3h4PntY5GViGR5pUSkdQSxkjM1galsPDy+qg
2/yyn89A8tHHaH0EGGJe5cPe89OiLKMQp1M2iETTGtz+JAwpk+87KdAj4OhLz7kPnEPPB4vGhbpw
6HuHfwuOZTYBw9I3b/C4cIzwzRooTpOB2RhqdfddVdEuMH6wf/kh8Z+MnKFU7YnJZc+cQ7An28na
FUVm59llfue9z4/6p3eIpStl79317Z4Is4TDJpX3uwRntITU6k0Gr4fhTJOxpd2T75tsM2s8lFA5
0f1dpn2b3Pt2HrHgF4sufLbsM4F1VRZEoG4C+Uxxmiwc3gsnhJr44Z4m/96CYR3C4/8wijChMIuT
0C8wASC6M/xwmMn7bZLEPopqVwi68kmWKQXWRD0525andr7XjRVtyLvVd9w0cYEuR6IRe2pAHiCz
xwV4YemXx9JFbsekl+nglnVQacY0Zxxpc778w+TlRaryH/iDO3H/vv5bNkdZ6I8P8+BuW4kfa8pf
bhiS2a1vDV6hAX0KsAhu7T4QqnlQbn20x0TmU2fE6R7JcJWv0ZRc/vlwJGavOijLZw2cjAXJNye2
znzxWHH5372n47NHCTQOJa93+RB/D2fO/kYqqMjEZsgLs8daI5k5+DtdEMfxCnH4QNqh0PCUfPZ7
b11nu7wxwKKaQJ4kalew8c9NA2BD7vNyfY2MnuaTGhI47lrvvaT0ipm4IWnSBqW6U6Ludo0TUZcF
lMcrjQhyMaopXW+n7IzfT+wDp1+fSk86Udfs+fraI5Lz1G6TFBjJcipLAzJbkJ0rrSPYOU7NRSWV
agm6FWQJIZbjIpq50tCkzZQDJ525bv9T0rS5MjcYpSLDRLFgL0Yf0/JJgZnS9T22T3E1FM/A11xy
3aznmr15ey+edyQ2Sj2DOM/4X5P4EqYHTV/dnI5tNBBgbD5MEHUDC4O3r2ualAruzwmxF04lX0wf
qO1MuiuLiFcoKZ3WlFqWNMK5jzh57NgGp2kWlEuw3j7BoZp+jMfjBhTVI9qof38cd+jKqL0dqNkR
pfseSex/P2zZxSYlCfIXYM2k+RyivE6xmOoEd924Qe6hv8eEZ5AWjGW2pRk60h/Y2tL9BViMVSRu
6yxSD8MrQVu8KHrAZ+AfNQjDxliej6vr0eIFwBCgZysWrEyAYAvS3HbxoB3ZnqBNDt1YQyZE/fFR
ty61Bk9bGv0N0rriJCcc47r005nl8yLaSRlEeBbvsOgWM9eF5/2vEQRFM/sGr33AQjXFTFfENIUh
iSldcU2SBCrCCIPYcIt+fUtJoZie6WjmUaDnNHaPmZ3nRPVHhqw9jRks/KYKN7ttr7jE7tUQTVC4
9pdPF9/5WuN2Mi8pThktyK+n742B24BWY7tO9OjE1tv2nTUtjWPgmBkPmNuJahNoBwjNEkVR8bDz
fx3ag1E5Dx0B+IKQ+JS5Su6I6KLKngn7oYZWdp5gMFfh/5MT97QXdBp82RzWXlER4fMzyYU5GBio
HdS5uJCrxUevf01sDEisJjBQxKJy2lxaeycmEUzEXS1vznLnxW796HaPaaUxqu6rm0T6wDwN/5PO
fOgJAo0zq/tBrSso1JHoalU3VRdALjuO3IcR2QyVb1xJlV0MfeHMEw3jnSPyQZL8uVj6EsMcfPVD
2pK1jRtI6YorA4oAYsYTky0giyKakgXcK7I7/LsHhieS/7gCumcRtScGYVV7Puc/klS+kZbkOKrb
8S8TnZiLbkjCdG+ud8VAGf23XHPI3V3HJbyS8YtvB6JRzucn6JM9IaOgXztJtVDGlKenTtVoxgvI
1XQO3CJOnUPStbNDBFv0UIjLZ5vniBtwK7z4Y1jxev2aAGXfhkmDuVgPelgTVIDL0SwyECRQyyE+
3Ngk+hcNJAmLGT0Q9s3Px850TUrtWGD8G+aLDPBnFKmYMJBxUHRjPj61HpSYbCZTMnDTpVbU+rZw
AvrthweIwHD0wm8+cfz2WtVUr5RVFuD5Cq0mTjmSLfibsfMb6W+OmPfGh0fF031s2ae3rfW7+56B
bvgDaCJQxwCLpjA0xWOaG7vU4bWYhteHO0gUaYD9b/Nydy1vWB0mO2ExIV3phCMV5Ibh5Tf7ckJ9
8gNHhZqXIBSUQZEDtbMC5ZnCxNxR8Qcj+29QT3p0zWVGUgFjxBMiHqvquJx9C0aAs1AjROm+FU0h
vOqj+uFNkMDHd47LNRtVg1Zd3eHMP1E1Ff9J9h+5oPqIT7wlKkSpUTzre/H3izqzWPruGSlwnJ8S
HglkHP0AI8/BY6VIKv3ycRZ6OGf/1i+VmEXBsqQswydAt+CLWt+A+eH6jDymn4gcMimoB5J4ngNz
sBCMKq+cBtc3/LY5u4arF1Y2Kg9iR4YdMrIzVtYbOSF43dkjE9+giQzX17DojUeigLSi9T4d27ca
jTHc21kwypjnPSusOy1zpqtLeqmq9vIPQ1FR4Ivh+T4kIy5LGfpAWcGQ3ZAUhJ36Kh6DkJEnGW1d
7XrpFO8BcdxfSQDQrfxy761orRChqMD2GZvqh7P8W54e12It3ybIpLusPd1TjFTvs3LzPEpJEzc0
xnUknJVxeF+RgmnrYvIxa/Gcp/aHkVXinVGK2bpOZPSv3EeSxfZc5BAm2P5ovVEBxKHQDuxfubeS
+l8yukvqRQvTZg9YWsa9Rg9UT1y2OccWs4O8wrPWoTyJ5viMf0D9UkDWZiKN7PvaE4Lsuc1V2YVV
CaP/HBuKXS/WZZs5VxWvLYnmgcsfMw277EFt0+VtqCiDVU0VCRQyWZWPlQ3V5rkXIyvm321AIVni
CNfSf75KvAiYfnXo8PDMWTzjP1jd4hgKwlXbbo5GABxdCLmTw2onPnEWJpIB5j87tdmz1DIZNqUG
PT/QwPkQr8V4Yd3Gmmb7aMCrjjaoIVYFzaattHC9F96xfofSjM6eQ3gB6TAl7CC996T31EYAlufq
PaZnT1pzf8OPtfpzrxZPLzF7/1gK/sdv9Hhx9ELgEOOwy1cGceNAuwbB1HSkWsCBNu34a4a24d2m
3tbrEDsOFyKoLevDRQihtZcwdgfUxuRHg2rtYIZl728vNxIJXD/p+29AR9FvqImVqBhsP3+GN2KH
42UmdTgVIAgw5LxZxD9mhOxrusA7Iy6XZyksjXc/qpjbHMdnuHhRLCLwxzCf8ud5kbj6Sov+Y0e+
oTPbxFyNGMBxsvQA0ZPLDWu+n6IxHVOxrF8dCqyIeXBZAtzA8JJXJZwBxwPE7R7/7C2zGp+PkvZO
GGcR1VoJ4JB5fCmp8Bn0e/IgShlfe1zcWjUKgxyXW69YD5RrxVPs/s7TP018u/PHn3hsDf8dXtrL
lQisULA7j7j5Gt9DQMng66JpG9T9Bb4h2jwnph69bbpXtiPmheT8xJZhamg+qSi1UIus39hBDtNQ
sObo99jiWig/1VnRwcXFKhomqtAUjHKAvTMLV1k4tDPycIeCYwWpScEoIpxtQhbgshicxeEzHxcZ
WEuUKytvS/8QcT6tcIYDj8NYWhXY0XLlyrNCGSmWig8HCz5+eYd9PxjxTrqjUrtEES669hEfXt0H
d/G+i1MhVtTyrndy23D6TiSt+i+nMJKF+o4uJuZlLPKEEqmX/k3L7yoPGefp6lqNb3Fk6dXftij1
g5XxVqWL9hC/qaIRO3UKJ5GACs4wD7uiKlKcnznMACqKVUU0kUfgyvr4vUUmeXDPA8ruPeQsxIy8
RfJ9tPYB/9ciCXhJGSoc8r3Do7h+O0QxFDtf9ppRKfeVsms4zcqb/1Cj4J9VghtZKFjaKQgdPHJM
5OSJIuwv+AWqATpHN8qQi81y3kGY2RxCp9kkWNeaRvlpQ5W0TgNLXkmbzH9emPymPT/aRe14IpVk
5ZSI08/bk6lGwqBtkB4ZR2XKMN8NW7v5pezmLt5uI3tks3fN0jxtMM6ErZHTnycRIcN1wm02Djqf
qB9mVtyycgq1EJ6f8Z+2Y35XKOiFA1Miwfdri3FTE9KG4Y7cwz0HDWn/zunUfHRloBgjU5LtyN29
A+gQn5HyYwtAOTfs1ER4o4B3xC6dP6P/KJZxdQhnqbP4uzwdWtBru7oHVS56wMIEAjYP/Ek5PXy6
vG9oA9q1GvTH9vPRqil9qZHcs1WHh8azhTngwgi4oIJ+mnzP9VGiaBCMoHdBJ3BunqpdaACaesEV
RRzGWxCJnZ3xL3r0jcM/t7FvnknHXAJw6ePNl7GHW+jL4FnBSw9iJTvuPGEibfnUTTx3yFDznA7R
Qshkgn6SDfavXhgElSrTGtQlC0FTHJxpE8wq0xNkHVJLLMsO7Z+7CFo3QRfNnrsoqZmvm8W/dpUn
MC8p8pO1XLxhph/9QB1Q4JFCBauAaxkZG3xcOahIyVPuk/mnWhEhjmUYrm0wfpCUmJKVK8+kCbYA
IQOzf3MjA9aoRbss+3rP5ne/KYpIBQ9kfmyDzVvs+SPzh7V7Jb4vZVE/8hrW8fy0R/9rT4SxVQ/q
ueXuKFt9lir3w0bEYswIBlsGJFZu0xw6EnTzMSvRU7UamY5ObijzE4ILmxrtATweg35ZNdh4BIVr
yPA8GzN5efWSRBs89ACUYrsxh/9CTtnjQaGy0s5jnYD7grt5r/u5NNLly4/m8AeBO/IGdzEPsSpA
ZSo3RYD/Fdqpv6OrwYhZlgqnjhXgsX+mLa4M06kFSeRr/bvNTWfkqeWUqbVnkTTcao99ufMpB4h0
89k2KPw/f0h63X2h+dvk7B7A4N7qMCmAESjaGT28+L/FCf2zrZAKND1D0i5wQgVR8x13k8MMsIwc
dul23SJ8mJxIrkGCts2lFHFwWnP9RFYDuKlkCGE8n3ve6F9LJtmtYtaJCapmPqN1Xhu5eeRG1tDO
tjXaHAInJwKVDL+k2QTk8rR2/8W6ee9I46nXlw5/tv4LRu68q2fTaMd5nWllvk/g7NttkEcoslAO
yZ8ZY48r9gdgmX2ex5+CceI9u0fr6UZs73UctyT4pruI8kgnvfkR4RL5+rjUwYKb11dcLnE/0AVi
FQJJ9eozJDzESB/WYvwwdNekJG6WKaq2GZA/+SV/XZDDzp7rhe2adNAgfbWk3/u3C/lBf9kvOwD0
2tLdkUYZm2seKtVvjwhpCZt/uPJR6hsvPXyg/lYQYiKJOs3CzOxYhvTnvDshhyeKanez53E4i4/B
IbKq+6HPY6+CXP4LuCbQi1dhbaerKZMEcpT8L2Cajqcj7v70uOGueHdoltHX+sroPTgj55AEDliI
G74goiKTqKdZtEZLR04XtTojmYiLwwEUsiRWvU31XuIWdEcR3I3thhgGpzvpNjZjTN71lpjN8rl2
vBu/lvsCAii0ollV6Pm9DNA/4CIiRXN2uFOd6vXq9fWQzrM944I2WMK+pH52jUz4v0fN51Hmcxug
MbqF059pWbdDdyT7y92NpJBlQeRkTLM9QBBd5sAJY8dcE8J47lIl0QXMysd50euWP9Q2tkrumTP2
XVFfsVGMOr1y5WJV8bMdMR3t7bt6yMpU+N4TJvQ1ABZTmMyT0+tX2uvUt6herWN6xfjON1lL5fw1
qTfrQ4PTw/x4WDAUoo2J7z0DoMBabOL0Q+OHu21TxeqD0uxeXg7OMvnWHcV6Zkyrmg4FnsPgP5XM
hk9Gk0bss3WG5+TMS9wJq7O1o1QEJ1E5MgZkGcAVCooHF1s5ozvRC0WJMQVNNHK/LJn1Iw3YvJvX
j84o7EaP9CS336Dkh/4t3z25hxGPG+K4f+/u//fZ5g5s77qM4T8cN3lW3cQyNE2nwFjmmqb+kll6
Y3DFHZTiQEonvh+pwn4yPjTvUTmuMZCVX8NdoTCF+ZslQ9o1kvCGYxQMGHbQmsYROGZgDVg270Rp
F5iDkqHANTsGT+Y2Gu7x4cdftD+5fGthK+ItRa7X2OsKohLIC8qIfJMHMxj4vxDUL1qFiIfnS9Zr
TKl9dGCFsn4tClgFF7bPCdhGpnvyD4EqBT4nV8zycR216KouN7bj8UGj8uFSUZe8jZ+qdP7GidkX
cmjjgW5cmM/dmwlG58lRQyjmmeUu09YODOlli2fQbF1MhNUJqctlRyVsmo5Yh96VCEZi0sgjMkWI
LiKLlmWgnV+3smbJWsG3+RY1wNv/MMGxVGgNTCDt4HhWlJX+gscl29FQ1E8rl52ADHiacVI7hIPr
mSXMrkTArKcPngxxZwnS9t6LJi/F0P2N6cTE/JRV9btjCZcQQxB+UKoQt7vaxbUHtZ2NCKNSjgZB
J0Vl9HLsAvmWdqL6kHIFK59HGHKzDYVTXNF0o4Vylxv4QUi/m4+O/nTSBGWVF1JvmAhyl6qof34B
UpaERhbuAKuVgZjiJUN0wqRX6+i7rS8NniA9lbytfklfRt8+ASTRzgLzhHSOB2wdRctbJl2/kuiC
a5QoVtHAKdTnkI4WkzOv+JGBnXI8w7SvbckqUS5nleNX69wA88r8bC/KRSuSVBkHKbjz5psvAAd8
GyiYbeiKZs15fH6IVY/lOQCniUJKuDxAUwuf4Y/JCafIDEY7lQD/M8rB5rMn7h7XWCq18qPORIZ/
PGClzzDIT4KNAuAU8pu00Zmtav9JGOYqQB+zwxMdlvojdIWAXAHmRTPuiMMCr+2gIytCpaM0HTVs
Rvo6KTLK6z6uee9lNULZIO8QvscXZbGz7K3iMSuVVxravMk2KbKczzyiq9v/S/1k5WKmB5LmgsKF
hWeWxIiOkrH6bsKjTcDRlwWmZm3HNQqBk+MobcCnx/bFnXKG+sz8TGG56OuSdt5/MD5z94HjiV8C
y9qDrY4PysNmPi5fhwnOVJbhbSYsXpNOyo5NhMETogXkHLQJ+QHha2VcVv8Isn3E1kljfYNqNGvx
xEGc5Yh0oBIXaTTvmT+LSP9pqBGfvVfLafD2cKtp3GaQfn9EVzT26rQoWVZXnQqcTGxR8lHoyfbE
QWzDK3QExwC7U9cYhXp3kt0uWAT8nnn5ZKcK6cOjHVB/vBHOf3l+1vKLiifvkUdK8HbO2WuTSomb
D3aSE1qFUT5ws4PwdoJw23yQOrnElAaw+vZOv+lwos1WrOD4vha2ahIFsoQfwDqwF9+3fJbRUGO9
ZKF60/omAhrgglgviltOegyy+LUo/9chMTTvVl4FRvjqHHxzIdI67aABOBOwRZZXoXWdRjwU24W9
wKJukdzIoFTLaCt6uPtcFP1wepCwpyNqpXWhZ70x0gkIxCXK6JeiJgSrrrSHuKeavl8v0azmH+3M
ct/LbmzdTENWiAMtcJkl1rASjmIiB83y++xltGm+EmIzEFOSJDIsJxj8NsJcnXaDP7N4KoopWEhn
B/+q5Zjs5ZcfI8mM2+uJcv2DKm+X144dn0AXgcfAczAItcjZjR0LKPFj0FG7WslvNBgWCoZL/51J
+v9LOyOq5aTos6ZD8e689EZ4XlPhu9/Ca3PEo9Yh8LF6JMJzDBIcPM0mdRwfZ8UY/TyoiE2K1CSO
XOfkHHcwQap5xJC53m8vFs8Y0fRePn1G/1BLZL5l9a2ESGZaGjF4lD5lFQJaNCCYx13locbG7GgN
wvt3FN9XDDrGsxX7yjVqJyGULkiOQxYfJDAX/y2+Bso3B0e6j7hZcvxieHFAjtkBgmTZ4qnMWGnR
tGEC/jq1FFzsdYGX5aW5M6SUDHUhhmTp4TEEBGjRo7rxGv09N/xNgEH+BY/IXuR/NZc0Og8b9vJ3
QHcGbpQk/9Earf1DR4mkBiTO3qQKoTKEvw4H5Y4P20VkIs/AFvOH3KS2t26dJmDqEj6UWvuVjt94
AamLFRiIC/ywK7Sj/dVJ+MLOuQ/dyzjM971POh9rPXcXvA9/lZZPlB0t2KXaPBoOdXc6JIKU6FDS
8subB9Ke4+Mj1htYePG2jF09FSD5a1T8KdPQ2tGcHW9M94fptM+cL+RM/UgpXqazV7vS0YYl1O1w
DjXdiJTV5lS/GQnGbDDGT1S15EJgkP4BD36mP/xP7YzaNaXz4xa5sj7Pw29UDXgL1P0bKAazlupU
vfPsCDVl2x/qjfIs/rb0LBwsyym1vqmFB5ogYg6GC4dDrjuhR13uCuS0M+elCvRQZB/wmLqT5tsQ
aPPg7ZylYNY0JI80tr8MY0gDGMyiGxkUWQQn5ipGYLbWbOf7vjcSntEprlBjbdFIKmw+PLd8LeE4
KKWHP60QAC7yeg44UIY4GAdGRSDfGt+GdL01eJ3/T3ltqfze4isUzPkC45MGgNckIscQi1GcYaVH
mnVogMbQi1HKQBAAcHSjUUOu4qpOqPm6QyBTTPwp27a7pGXF4mVkVfTSfVSqyTEN8svRmB+zBYvN
kzTWjyZASUIsA1jyPlPi88WJDcdl5rke7AB9QSbuml8QJG6wloK7TzwmfMvtHYEO5hYU97gYGBlZ
NlSbM55UqinKcnZ+CnareOXZ4G6RviqLwv74ehuQwcwmCpJy/sZVIkyGZ7nKImgdyFvOh58LTMFB
riZEGKNKJuw96RdGjmQ1M+xge/svZ4G6wJAZJqij9y0z4qIj/xVs4YPLutWxnEMPg3idgvLF83mT
g+x2EWDC9CM2hNekJV/fHKgzen6gUKHPRjKYppaiiub72WJJOAR/TGocxJE8uGyWrA32BxYiKE+P
WJJNHx8qhvmJsQJ/RswD7WNfFiP4XIwH/JUqvdXB9H9/q1WOa34fQZPBuqXXAoRQSEvjHBtqpb/i
724eddNMGHzc+07P7iGicVpt/jClYqYy92xKlf0fFUe6RtStH3YZy4SpgEJg/L3XCh2VbFeJbm63
LJT0wAgbgoa+nCcD8ZCVZhYPQeKR21gMh5334hkUolzxd/ygdZtA/KNrhNoH3Jz1zif/tiSlEAOh
WfjW3ogo+/o8vJREMwEUaB7b6Yi/8V4jY8q/1EAjpTZN6Kg+NoPvQiY4lekRaciKxx7Wk8nM6srL
SzaBXQUiPyWuJe7S4Pol50gCOr5mE+CQ7qRh5DWZj5O5HcMgct7298IhciY7eSODaH8JLxVvv5M7
AIsWUsh6I+LuPpOHuxSHuiQU8NMMAJO1o5QENaR1gCX2avCojVrk3GfRNot0wt9FYtF2O8TV9+Uu
873Vl0vvS3J753jALbS9SIQRKBBXpIuW4ElfregOqBnalFwNy9XMA7MDRrQ5guLY2IzX8/bxNfCG
y11+6JxY2PseOEMkC4PRvtFG7ANJjq7xSPRzSiQpij5ZHK7Rn3UZYFdcRrk0qjapsS9OLXHMRgAf
wsYQQ5H7GcPu78s7laHN9PzHtERERcc41ntOzVYCC86bmWoppLC5PvulDfZnRE3MJirw3Nop8JzR
VOt2FgxUVcx0wG1NrNkebhVROtliTGhkvp5i+CSxRHFj7mdVJTldI1nQ9AHP5kDVcEVIcZHe+YYn
tUzzUt6rCKdk0vD7sTq5OQqoUUmPy2/X3OAMeup3FUJ5LqClmyROwuEcau2L4+EnzxCh4d+4YuM+
dmDOrdMCTtppGbXW1mUry8tR2Xz69ZvdoBXP6VvKBTv5jl6laQfPbuD2FsteLi2lfAT2+mw2Kg7J
iWYQ54+E2f36Qbfwjd/886U2mqszCZZhqFnSdLnQIw8r9WlcZoK9egSRNRMFetPGQZoo5zia6pH6
dXxeZectiBhsk3EpDzT00E8KmUPHhIgD9rAzVj2noVvs8ceBgty2ZHqYVkSltAAHoJbbw6lu5W2m
LewAumMCpR9poJbUMG5nRniAcgpchqWkxOERsvVzm5jHEq6EPBXie13TPxSO7yyhhSlWb71e8VBX
PCSbWExhX9qbNyFlINCOJQchbTW/ClTrrCkw2GiGeIX2EV3JSXmIuI/Byz5nb3XJf6EL3WyRDJMY
t6sZcDDrl1Q+xiqd/qB1gbE1TUPP1M5a/MbTkp1YMWwQwuWh7zPyeskN1MMAkrn2+kGOaTS69o4L
oq/6YTgSJItQ5WHv50G8/CKkZOG6KD3MO4Ntl4Gpp9d+yMs24BHOywdVUjGXYaeM50G0t44eTogf
nBu0rlvAZ8gZTdO4HuOtzXUIEraCiEV3a6jZbayOKLZojS0ABTQLysXeiom52secTOCsc6XoGVAl
PM/ymq0RCTozjGsK9fRhHrC+jr9W4n9zjWs3OmpDuvNHRcMLUYo+rdiwznquP5m+dqe5jmUGA0Xz
Myg5Zc8OZ05gErKUty5BsknyWkfcFLPnuJOgufMq2YX8gKZY5DKbplxk6oKNuWahuQB6sudZVipO
HZkTSqy6Syx4iMGeEhhlPPbNyZFgsneozH/v0aIOVLiE3PwDL8HFS3ge1g3ltxz6visvhXOdFGVE
/E8dTV8+kvZJyrhqiE3N7uPr5afYjxvMHwCzw//3a6lPPN9cd+stQLsym1SdMCoAC2efRYWro/R+
Y98KqgzM6BxlgJ/SgFVPyU/X+p/xdSK8YfirlNGHi1tXesalXOoa9m9MdiF12HLfUchBoHQn9qZJ
VMJlmg7mbK2QmRUKAmiMpTTKIfZdhntrb8Qu2Ay28B3v/zpvTAu++sFldW6boZrV48vqM+JY+XWQ
kiweN+DGcVaYZF9rABX+yUUZ2rqjFMiJ1063mzmL9K3XGGyuybLHoIcLJ6IWF5DkpWFRCYPpRFts
hNYOb31Zukz1RauXnByW4PVmzY9SgJg+fj03/m6HGjkyUjR/MKLe3gg3wLtnxu3mykN8fs9+2kLj
Ow2JIZSRL1sGaNy3VvZcQLMgpYaD+npRGPfeksa/siVoGw3E0jVWfHz0OjFjfJhWso3BnA6KayXI
5Dh1StWj6XYeQsui6PNVfXXxLbBB64pouPELUXwZLMmCEMvE1e7FTbQiR0Nb11Ngo5bm+36oMK45
GZt50wgqz81QZlchEZA1PTzd0CF93WGhNAnBCF3dDXbyH3HHZoBJSH6h89aN0dEYMrq1u04JgpXL
Io5A+MuZLuId9aF9Eu32o4Oc2lavenP6/VR1JoYXvg0NNBhpUktADW6lzF3CtluhrVDOao6LFC73
OupEwzzUIdHz09rzcWlIZ7rs4QhwHNtZq+XqzBoxj5PBIv1Tv4bC0KUw6DPmRdVh1g03C0rG3cZU
+E1K0161YgDtST1mF2dvq4r4USAe2/FPgqpjy8yYamOpJG/G2XINYLp7KIy3QVeh3WKsolowXLfI
ohcCUB1lc0S5VTGxrG8CoQjgeRjfl9OmY/S9USVNJ472Nq9pFkZ36u05PmwS6IFmyw5JcTTQvTSE
nYyNSOHyUKskJVa/X0FECBwq0Mn+5e2mmXV/L9FBeUb0U5CR6H0wIS6IOjA6icQAhTQMszT3TJ3P
PtA6h09JqMUeq2aWHw/Uir3vVeMFkk+UY3Ecewhz+xwL5JLiF1TLjygZsTEdF0bymWNFX+VLvDcI
sEmrcuvFauPEWO+cJCE+gEm9Cm0LrVMwIjWjFEXnMPDjAJwB+Xm403rXjwFst9bXml03p2i2CWH3
Zmdzh1sv9XDu2J1aAmlXgCzuHhpDSfT8NISwymVHEAb4pdLLl/4JMitPeY+B7t1JcomCrv9s0Bwv
no/THXXWQm4y8oAhKdjPEUJIRIhH7MxPvJzQJJ7AIbZweHdGg/Am9snSEYjTNN5GYOuocwvRMIej
PLYWvYlYUpxC7fvhjP1qwCulKCIW7G7J1LIe34qOtkUoe722Y9oILDWH2DzOmn9Tw8V8FASs6P/+
9hsHLR/tIUvU8nkqGg4QwIbDMOoe82HbjABv8CqviGL1Z8rD8ZOM3S/eibGFm1wQEN9WqDtml2jI
aHLkt6BbYn4qIB7L6T6Ryeyygp4mgK+QwNVMWNYNRnIVRKmd+1GleR2eGrgqZ4SaU0OLdrblohhL
EAYvDX5fEox10zc8uEQqfOpZD0ds/+3K5qziZdEJpRWTSOkOYLzK7d8UnwRS2bq61OsxSIKf/hFa
RfG0eBVD3bQhs0b6WrUS+NgNOsCuu31hCu+Rv13OUifCRsGHASuAo4UE+Up5ANfEYFNs2sIuzoW3
bo5kH8J48vUiz3ovwg2WnpnkeS9DS1kZMj/s2yMYEshZxT016zDIU6IzLPrz3NYe4LCBLFUbI0gr
OyraXBCB9S/Nbn/ffXtWck6DDaWepVPYikbCK27RSeC3YxVZc3yAk3JaEuEwUd5ILSGumUWO/EEr
7p0iv3se8/Lg+Lm6wt2nSC/qO6nvZoLZN01PUacbTVgmMb8rY8FWN9bD8qF8et5WqEf6gbW+njNP
MjBqNN6/2ZC/Sk4FmTxQ+oXPO0BNpy2amrCaLeyzi5GOR3gs2iXGqr7XYLHiOGxiqbst11sf6jPV
Bg2ugzDY+9BDW61rE4KQE7x36jKdZQnHRtB1CsCGpMPFhr3+8Rboa3jymZJZzUPO/9CghWfT4vkE
EyuyDb+qDmbj8zeZt6qi1KCM9YEPv+1LXoO4kpqsObajOw1+1KgJ3okH/y9ysHB6Pr0jqYP9X18q
Qo/57bIcxR0bCPotu3AE3Dq7ypT0Tb4L2p67MHku9SuO8OvvT6/yHhypzt3jXF1BwQFwtMi02ylt
W1BBuJVVbuSmMiFt7hoRyJQv9liyzFrfeFIUQpEB9JeTwk5e5sPJDBsn9zEGHBWxe3BlYcZKUTtQ
Yr/DobNDZJBmct8Hk6ljuVXbCMyqIdtul5cQZFZe+nDsXgRMsmkOkZy/UdSNBP2F+/6l6BpYpwZ4
sEF0gRPz30KZSx0FUPcd7/wsy70WS6ktnREkF5Rkd7r6nH9mjbgDVVuH0gmLete7b8NFcE+U07Ae
ZnXTYkxiYXzYzCEu486F82DzXdb2NIqJJo0jAkvpWj/tavW8VUMzzYJ3HBWh3+gf2teNU8PrNP6i
BOTUt7ToZ+npDAqQp+TfAhYWj2BXL6F5EmDdsmY0/JlMVbEkUDgyIXiziALpuDrWL6J6ibeLpdaW
8YeFPIz/WyZ0/oKy5gFFiVDS91InTqQtOtMpGyJM8YuGdsRgZZskvbQtqGqZ+h09DSqcFQlnpS1b
LMLA7gPO9qDKHppG839u3CBBEbmCHMBnhN1MD2unpm7Fkt1nLnnSGHd5Q4s9RjIcU8H7w078eZIy
WmvolPlPNCt3DYSY8m0sVJGZe5k63g6iFN25p+0+3sJ1by2Y5/5F2zjfH+J/KFLJ3xAtaYQoLLd6
Sv0BquxFkSTCLcIRurCbb5WExU9PC1qWO9Otcmc1HMVbwXGy3mVSD5qP5Ufo8Om1RaQZkh/2Wk0G
YiN5d715N1X0UingbVp0W163G7uNZn5GUqc6ro6gaqH26XFIgDR7JIjwmqMlwERnsVEbX1WweQl9
zTeKGlSeEENP2ADwHzRDA4uqTvpvSkiRnxdpHL0mlBMjprYScQ/cHEDxDtLGvfAyK+WkJF7EIfZg
1GAsQiNvXCfXyyTpXo0GMu+E3zymifLxDhdusNVLG1aWzt3Ukh5qaF+TsyBgRZuw+ta/akVCFFOv
lb3YmveFHgttRBatUzcDN99GtdFWHOy3ZzQYkhPDLYc22W/LJ7VEpsen8pDt4TkrTj4t3U9sj8vN
lU9ATG4IGkGoDN2ut1wppiHvDdm38PQjLlJrsHyUE7SL9F69en9ajhf8acp7eTHsD8Ex9cNHXWA1
PCvmNM6IvRuhGnZMdnxhvhQx8bmr8sYGGVqCeWFY3r2GD2uDVB0PL6gTuT7WnhASC9bA5pTvccOo
/hy7+0FAE0OtwFOCLkDAiIU5tJQijK4rB+CntGgJiQWyMlOOyw0NXz6F3GOoO+ydPKynFnPdQuDj
1cSwW9PYViGchtbeEZHv5oMaDn5x3lyI6DJPHFM86jkTz2Ed/EVi+vCWZ1uf6D63IYyfO+yG6bMu
AfmiERtbsIzImE/kpnI5XL4RNUBl2pCLg1rY1CDjcJmGAyHb9QGY4ul3qZaWNSIccoDjH4nK/UjR
+MGYu5e9fCdyYFNmaToER+8caSnhd3xvpPh/VoWchyM2/ANIyFmfdAWPhdgZ36cCjXCYP6wPaSij
ROC9sXe1jBsw1dy5WbprSimU8RPVl3YlFPvSts3bL51wr8wNfUMQwSqOIUdbWxoSCwK4E7WdAFDF
VccFu3tiFkykjzmszxOAjeEktUo8+6zQiWulxmdUJWfqXBFG0OKh6uEzqoGjVwUntH2mlvSvSDmA
PvuttLbKid5EHAMWmJYO/K6ALYuvLZIj12vLtXuqDoqnD7+oUt5sJGrFD+GP7fboaZsn44lPSgoH
+g/w130IXE4dmT3fn7rcVOfE848CVup9eBLMOIhXahMN7RJn4KphiRQ/XmPtA9PgJoBxfOD0A8io
5idN2gV5pZ/b4/KjLbhUCG4FohpKdS0jMAGj65ZdGxlZC7hGVvFGo2fjC3Wkp0jIjAhd3HV8PZG8
5VxyVzaXLq5xn6bAWHgKPsyngrrwNmubOpF7gDUpPXTZ2R6EOsUoiMLZhDOTTD+caxBjGXcnVInn
njF48Su7vm+DfaIKtdD6P28GSsVUi0Ql3/IvUg2gZRJNMaGx2kSVCKBO5FfB7uWszVKacJgmn92a
jMtRTRXlkuvtN0r2jgqD/zD+uYoH8eJdlyXWv9v5r3f+DXN7eDLX0UX1N04P51fOl9bBnK3JwhHh
WHA/7tAlrBpHt0P+QNwqNBY0Oul8v5utgaDwx0DzX7hkhxwy30jzOyENjpp12FNsLmlIhGoNZm1F
K/b8i/iuy1ntvc3SDHI6NiI4YpgzVqktrjgQlGadRnGknCbyEWRsZBIyvoC87SzaWNalGjz8FX9M
qyl516+FuKMF7mT5dUBdRciafo1uMHYPeP3l5fo6lBGN3V/JPwgUSPk+TF2QhPSMbsDhhnKdFrKG
KZuyTVP+Ktvxb7LBoBB8TGJ0g7tjjpnbkZWqylrvA3kgPLiifnWYD9ezblxJl7aoE/EwqcI2P/5m
Hc06tgzuaU7lKuQ9tB4KgXnfYr275E98WcS8Mm69//ZhxoCK48vJ15hAT5EtdOj0VwR2Ys+UIhvl
TJFhN0hHMsyqszfxTQeJfQKcd3SpJQWEPtAKdDhEbGtPWLsuG79Wfjr8XJQ2VY90DGXUYXusJyEi
RWiRomikOuBGatCQo3P87wBtDWSsk/7b2H2edDl5X9cgphd82mnu5fADZztT9Sc4PSIenk0XT4st
ZgMsSnMdHt8yuqec4Ef3Vl2BeAQQREFDE585pO8swW2nTjScJMKQMuX+SzrTPsfkOahjUd5vj3ha
FEBmtuBEkivzFznBZZzJvQx+2+K+jYpxwqAOjpdsxmcAP/wbFFzcNSpu9tdnuf2PaWMI6WiCR7l1
ew23MWnx1XZT5BoaWtUkt+Y50I7X7d+CWEkuj6l3ljpYaAGObcyI7D4/2nF4kbud6O43l/UGDHLt
Lpin28gLKNNUdXX0anviJ6Eh7FLk33FAHYrvBYEFtyV5Jv7gCPMvmm73nuGD1kS63odUtSOdCXxs
AYtHAhqvuRc2UhHz7B4hGD/yDE2mzDbtByHSaN5tNwoqVh4v5tqJgGzN5qLKNBw4x8P/U1Ho33W5
wPVJrfY6agH38OvjgQr/H0tnkg9Z7cHZvHBVM9tGZYGbg1hMcW+Q16Q9AvS9oDELIqKzy2aT3kRA
3hWNjMgT4xoOAf8N8Q+2lF8k5WiwyXx3/r5eBThPufhA379WDpx8QlsHdXl0fpLyGHCiwPLvIO7O
r3YSyyEzbXQodnN8mRzoh39P0zkmVgr/H+qbjJhA3znESgzXV4ONSsdpC6nzjqxCV5Pi+IXbftOw
70C/k/D3gfv5EgLGWr5DbyS+60UwfMtDldAjaEtCbWEGFXOS2dhiG5Q+4O30YLV/xJtE/1eGg63u
BdPgjgdbi1+lBnZUkb6mzERYOodSLQnVGz77eyzg3E9OTGqI2DcZSM/1bQWJzw7mI7ralF3QnPGN
5R95S0Y127vD+qLlEY0VyPNPx6J3MivoEXpIHRPuLYD9LJvO2LcE/TayP1pyrvFmtSHvFEpvk8PO
hQOWhk2hJ+Ka82+Tw9gtdZ73d3vIEGEpixw97NT7uYzhHFSqBqrYap8B/qcpPYtfmn7KRDrHwqII
ODRjxTeQp+w3GWi4LdYvsIKXzXhmETDAPWbSXqZadeUdiTBlzywFgNislkxg0fbHKY5N0Bwy3zZ6
bsc8TY7/7aQLUVKJmm4IB/MrUijMNHT3jLsj5zW11c3GlmHimT67ki6Olr3UZ4z/1ufDv8IciMP4
wwbgGEjxMbemkTDQw94HHnQqGIIC9/YqiDVXnSQ49BP/a+ue5EJvFUgZuuCIGq1Z+LBfUOOPN2kg
/s2SqsnZdPj5xofp7L1mJxpXy67xTJUoYtUYp9Drq3QuZhPCbyeZN/8gA3vObv3sa+evy8FJX6wd
tRxDydnj0lUimvf6o+bcS99Wj1ZRJQS/V1Cwwz2+uQewjq9sY71nFukHQU+1KvULsq5kPRBigtsb
ddiYIXN4Ca9bTtpk2bXIZV8oDDOLh9zCMbJceG9ix0t8Bt+EqczHUPWIUhdN0d0hhLVjUZ6uQ8F9
2dhaaR+iHWkiWJlLjdBxZiGUnxLMdDHiUsFyMtu7RZNdN9WHwARWWOR5dcWtv49RHnIswxLKtRie
iJ4KLAK0wZaehRCvJ77Byi51UV3cBNKdEMlPrVtwPvamacyKfyHXowAWoJjp09AiN+Lm8ElTyO/J
aJ9bPcfvvRn374lrQnXioU1KT5+yhMT0m9DwwnmUYCC69rfYfJxyAnY/irLep1QLdprN5DTvcV1c
OGmZbpDTR/Q/IEsSgD7qpuNM2bgu8JG+zuINdnoL1QvgGkSkVtnz5pHY+2+wUgskAIggcSRiRMU5
qCsYtuB1DZIcca0hpfj2dmxXnVQY5GTgldzjkl8J4c2rMdyyQwXE0HCfKvZuk1kyfSFXtP2ZLDiz
man7St2L8YUcs8ZSJlOzKMqLPVghhcnwzMmrz6EzGdXLfIaY8g3WqACpnzlEiXXLwWeUDOA1Vz3F
dtX5nGFSrSdKULHtSrPfJAnKNvJ7EZnZrJEUEhUvHMK6XuUykQG42mlt+ML6KEuvQeB1eX4tedTd
ySNTYwOZI86/kIR30EC36XbbssuP6yVBCXtjnTsDkbfPuS93O1eot+JtMmorCXgEL9G/To9Rl3QU
Ah4n9sbnoEpiuBJXpYofWQKSDWWL5TsO8AjvacBcw3h+5SNVUaDHmrn76A65puLzV3dE8Pbz6QWX
PBiqT5l1vJy4U7zEQA9eOc0c52i7Oxo0JLFUGAfN4mc8dWOQob+UJXZlMez2pKXOKpw8lx0XRg3o
QIqq8X8R8/GWvvMlDCn9f28o++gR+pCXLy0VPloFHRhPy6fEo2v7WMv+Vxi1eI/hjVrKKqk5aUA0
518A0MubJJM7LR5iGfenFIqoFqf7Zeq+pd9qW9+OsUXG6UKSCWF65hMONHBJYFjmxSwi27aOZwT2
w9AaPeIg51Il5qA8OYQCO2TmlDsE6uQL//pSAebw+AFpukidAz9EGbQnvimLCojDHC7XOizrfXgK
H5OPB/HLTemlzouMZ9pKF1rSy9zs4MTIFNBvWSt8tUzlyZtzxYXIlEybKzQQRlJpQaKaWv0suCjk
PlgISSlboHATwZaH+KfYtTR8VPhnvm/BHL/BqrRorYKDwl2F6yR2eWcLTiBiNAZ9AfPuVFadK4a/
Z1ghtWFGZgfNH0Z1C2MBI9yJA2GUleSJlzeyzzjfW375citi3FayCNTFKU6fqB2WueWywba61xfJ
OGgOwXusNKGlMq8jK5YjeqaApdhu0osSI8A/sdnytwnkfugVCMGZUJIQF5nkWFFJFXEN0xEDK3DM
+OEGdaHhlNv7t20IrySDJKHHdbMGjKwtWii3kaS6aeiZVB6CnXXuOYMhUiTG/2v0S+AC3EmEYjzr
hP2vanhYHGepbRlQwOZX2UA9RO/qwy6cXcpIxhxKDAORGs9kI37M9r+kf0uGT772+2UftNjmSPl+
DbJ3JixKSdFRLbiYrH5dGnN/VdEEb1tiHTjrR3nWvGaBUIOLCP+nMxxk0cPiyKANuOlG4hBJgt1C
q1dj67fx2Uo5DfIw882T99O7fzWGV/vbYtzjdzMgPvpM2Fb1AwNfG6FcWicRtVeJfhuEgBPeZeTL
cQBBs3XhtyPtMacPykDqPTKywEi1fMJgDTQAERGRPW8XsIigka579I5JOA+F+EwnKoDl2IUwmXHP
L/sZRPXw3o5txNKGQpkvMhHfd8/TyqkQKfolO9MFm8FmxqKtnAM9Bsz0k9qILuMDaYQryXAiPpE3
B25Z/jHozud8g+y05xsC2l2eCojKiP9YKPIW2vByOOtNeWcTg65tCkWZxE3POvoErWDt/uJ/2Vcs
2bgQcHkzHBEf64fPLT1nyoHHnTZrQK/GcfxQ+RJuzumPWOJVfk1an/XbXKG8EPYG2Ql9d8MCOyE6
sRveNTT7iplTgNDzrVBxXUNVKPJI3qtB1pD4hyzkJdHha78flITHpz28p7S3sIWJgmuz0L6KZrJy
ySACIVXstIi6ubkLUuKG9cW+sTnSpDga3RSNzX0SJXWFBnCVI4qr9hZDjDnIXvX5VAt3yZNXYZO1
Y4JZq2jaGRtBkC2555W/KPjo+7obByGvNqNdvJnqBefRMSFT3o25APqzWi3CSwHoD9jCp5Zjbwvj
0VuDfBnfqnCSQ7IY63nL4QnP1LWA25NFFn3+nP3+Oznx3rE51mrLIHDyF5su/ALm36neTc2Vta8t
dxhRAqZob/EvebWT0D9acVkbEKv9wKYrRQ8RiGD2oNwRoPMO1H1/W/Mon3Jo+sanoZAgStFO8zax
XKlxfwCE7w6GRGzYt8WoPnKRlIKJCGI22i1atYn5egpgLOa9NlhNwMoyW8906qHkGUj//r+r2MOP
cWhtszTL7n5atzc0ee2TcS3u5WyMx+swZg+38x1gv+Rle5c7VmMDy99qS0jP8SZvEEG+TrcWXMAa
s+N5h8fuXdT97tsDg9hhvxhc0Cr0D+T+eJUDg5Zqu8KoqyHja/S2D2Mm3X4e/NwJLUjGvPy2e/+L
Bp7OKsLfc6fCvbnYtfGBsndj0wz/0gtDCje0JNi53ASWZybLFUbgKYvN0tifpwqAhCW3y6MzARyU
Caiauxlmay2LtSjKdRyVB5xY3Yvn/9VPmXWGJH/eH4A6ro2BInfTy7YwkvUPtDUbxbwTVfaAZzoF
Xzju90FkV2B5vvHdF4KsvKcNG30KSJJALzBuYa5fWjfGRb1LO/FXKOvoVcI872OhQrZhVcsCAGg8
9r0PCxGiEEndPFndAbViHAOClTMf4RcNSfo/10X+vB/F4xT04ddcMJDpNC4XGgegvN4Rb2J7s0bn
gCHx7FXVs7i84O4w+Li/PJgmr+HP2T8GNdR6CcVmFnsCujl0QsehWpKJV3u3tb8ocpirzcJtKRSS
RBlAjUdL1ppMbMPPjQv76Q+tN92jQnCf/9Ez9EEzSKzc1PCZlzRQbn7xcgBMiaby8woumEHBk8TC
ceTEqOocddHH7pggjEaT0SuVtNvCf5FppxTEEGn41DI2SN8bVEyFmLwb1L7RyXoqHFa6SrAluTEw
OQc34Yj1Bs1zoNg2/m1C4zNxA2AbqDxUw7MPZo+ILckbDW2BkzXoj7Uca/nr4TVxkQYB8gxR27Xa
+katiycmmaHSpKsjaLGfAYgIRL0c36rkIRBT/znSi/u2ecNaj8p2oDGPiijconhsErrHk0YCDfRH
qZkeziPAIidbK3Hb/Umri9q1QIzbwhTTCevpfm5nx7Z2ez0mnGCQ4QoGkI041iCE4eZ3KQqelyzZ
6N50hLrHggqpaH+rIx2VR0RgOi2//3qIE5vbv6AqI8Jb5+lGvlTL+zN2Eq5LERJ++NHXSMCdyPvt
XsHgDegIefYyz1njPb/9QnmHldu6+2QoD4bU7bnEo100VBRLXLJSQ6PLNmv7NnpJt4mJBsGFX1a8
uMUIHK8pNeGA4Bn+hzVOp2ELyjoju7aVXMVrBzWVoQstbAYBy/x/LwdoQWvHCSfKpWCiTLmMgdJb
qioQ5rFxNgW6y4nTrmmj8NEzMV3rsS+AedP/RUdibaFoKnnihvsOkdlislaBLDybDPPYhEP8pCtN
vCu64ndssDH9dsLl1H++JDvxjxhf+YOViBzZsYARY1SX0wS9yiEFmmaPT3KJtf2zeLRCjjjCtu4u
RLmFjD8tHZd1rO4EU1Piu77d1qgapu+8frPWo/3ImKn0lTaZrjJ95dqmp1XRAWQZQouQMHGzE9Df
E5wfrKRq0qLOXGiuVYDUGDHi5cIvVmImD+A2OxryYZgskEI4q8GpJmA7cTGtZFJoyUZo2uEdm5t9
nbqijVvz9YOLQeQRtEP+oYYXn61x7XIOWSPYdeN4ehNLcGcZ/E70mpxbXaQ2ePg2UBme5a3R6u/e
HXAqRsVK3oT84VF4PSjqJsl11WTTbR8MlhgIVduqW/0af/V6w/vrenbKutfcrxX+b6S1CfehrLgQ
erkYY1B5ZfoemsMaotKr6aamjZcBr78yH8tt7p5Km7cdj1sOn7llPNiyaDoBjbE5sQNM3+ih8w0O
ApFLOzLC7aWeE/xVkLyq188bdgtviNYs+j/m5WNlVuB+uTxiqR0EvQNFKlXy0TqddxqOvHOWrCvT
yNrC14RnoN/cC6oaLKkDXYSnCYR7Ou/08MboH2y0NXxmZR65Ti01G8m0ORZAkFnFC6XMmzEUMgNu
GmRkxGTTsZstFPSmu8tSP2No96n1E4vSzPH9hh3j/erj0O6p2AYloJ8TrVKaxQJXB12HmWjYoAl9
w43pHeKfYMmXei+Ec8b5xsZarkAk9803vm+u/ok0HxSSS2S7JknauwZst135ISCc9w3k+Y8RWzsb
YXX9vwwylZZGcGF44/2/QVUDtFbF2IH1zZp8ISZNsFi3Qco866Fe7R0pS6b/zDzJgNGn2t5WJc7O
yRA36mxVkqHP6ItiiJtijOkMNWT5S2kyRj+K+FuwcdBauaE0WRESzyADtip+KuLKjuYQF8xPByyT
Zd2o51w3+GgrsMwVl/rcqg6i57ZCDJApD4aSHa+SL9RNYXURAYc1QRTFICVtNXIH/cJO00N/z3ab
4nN4Ij/Qqu9Gzrna7CO6fPbNzrQBsxwna64xEvDQyFYyLcaNNoL7EXCuG5YWcnD1cbITnILENHtk
bkBW9xqsummGWxnicUU7Q/Vm7IpliawfWtgSssQYGVivMLmkwhTfBug+1WUosWS9gS0flWntZCw3
n/3wov7ZuXSTnm2IDR7OHQ/51zU5FG2T5qaHciSgIPjVQbwl+PrsM3ozfaZcorDxQP+aKE8NUCZD
m+UY5+5IQz0Xb+fXx0u9CjQDzsVSdIVgIEJIBvyH+pIlwKRpAm/ybUSGIc2HUcRuI5XYHbjk0TQU
ZRmN0fFHAuypOkOna+cc93Nkw2fAY66B2ZpWP/uoGPCNEDrIPWwrHgTUtKh1m+fh3O0UxeNshiEZ
J6hgkN17iFFeLvtmqUGV3sHfZyMDRSPFp/+RfzX0Xi37zsPI/LgKACRXjfaSD7Egmq+FeBjQ8Xc5
HmxfMt/81q4Dzk3/x/KUr2z7cjKgWBHEe0jgtgepGxnkjcgt4vWcUGL17ANVuCSfwrI3di5I23Pa
+yOZEPqN/ElxCqCFqmCNKEPihJGEepjegOHtsmK1NPa1tqILlnK3NwDd3ZpYSZt2d0ezCPRIrvn3
nAiV7ZuHi8WaGaCf+v9JuT6AOFL7BW6tCTumyZLgxyJCjqq3/5DxV2FAtgDPTDifauB67KiFMzeW
WnYTLRVMAbsHITKYeT8+wv4hfBfF+uB9YzFC5E4BxtyJtHj0aNlO/7+pxfSGfPVm4yu3Q+Lo1qDO
DHY01Yc2lw+U+q67sfogkf3vHwv6mfkN2jB58A/4m4b1HozL72NoG9rU+IbRIPyg8SIyzLqNEo3b
r8umb6JcgITeCNjmKt/QrGya+bC4RCDtVwNkwf+dFb24o13FVIye8hvRjQuByTWIuMfb5KXYCUJF
zTRthcPQCJJw6IaH4UQO0cnaNhuS3+Snx/znqUgj/Q1zFP6lvd/KVq3oJD837u4B7HKgui532bo9
g0iX7osvKre/7GSDktt9J0W5eK009uGtej1H19xZL15DiyTW0AZo5QReYvVf7SZvc04QWO+ZJnmz
GslBR1gXY8KCWgq6yHN0z/rXsiKOubrtF/1tnq0TkSsl8I4M7bOV6Az15F42OCaGjJMn6AIk+GdS
GXQxsBI3oeZVVkMfwNI+Jc+RtybsHf2iCge7t30QC6PqBPv3PAUPq+TzLrwIZwyzs+aRJDBEmTp9
z/qoif0BDcp8mOV28HcWR+65XwwpYT/7R3+jqgl9+UZNPTZ/QN6+e4DYe2/9z8ACYdoNQ87RBYde
eChXL3KMqfYpg+DoOuH7KOTqMSiYYKqdjp+7rC4Cht4lIEsos1G5tz9Juo5bXC7wrq8VxBGxKfg4
nztrMijHgEV51mtlKHfmSaXA5D9QFk0AmehWfc647YP/SSY9QMsGqsZo6GQeDGJgr3cVw5AJZHwd
qGjIY4+E4aKSj2w1bn1Utifk8dVNqxgckbiclc4e0Yb+wJk1eFJejRKKpIzGw6N6RfAWtdj7SFf5
3xS0qTuBIG5Ol/dVd+FxgfQNiHSfgJgdjULcFSIT9rftWe3eQUF6W9Mj5/ostd20LM/bUE5v0xWu
YB4egeEOckvWfeh4rxq/bmHqGPyu6xt/etbogzoefhBEtWGIdbsYE3MflDViS2pfFl7DvRrsP/5q
U46YtMLpgRAi4eHbXPEXOy/0PiCDQyPG41UiVbdGiDLZpfpH0QQJHZ2IiWtHcYl6A16XiqtjFb61
627B7w/L/vrXUv45IGoxbQSACIjI7a92+x98RgMXEo/sYO1SFgIEDRIMmp+MvlvDhqofhD5UPoAl
vzXp0MlCCE215VzlGDYCiZH8isEFsJgTMzg85uy99gIk84GRd3FiJEAYOxMWOUsE7uLKQkFYtSl2
anCEt80FqO2drlQ5on40oAmEWmZdN7fiClg+UBKN8Yr4EABG1Iu33cycxFulozamVgTuywhgkPI9
myA3nAhpOBodWRkVazJlnc1pemPlZhjibPoQ9ST8P8fLGdpfvN/yWiyXfVTGVn8ptlD3j+/7C23n
C9AmiJgEG5URTd/FQ027TqZGHSNs35nU7shvZj5EZ9RAXf12FS0ffK8hxmiV3aBqmZzVK2RqxR5V
B7/TIdJ+3Uts64PAdf7WwMk6IUHDfFpWFdAcU0hlL8vWqGjvBygVupk47VPlu6iWF5l8FjT5Bxxk
UgwY34E9JHqML8Xv7hlou9NYerFVGNB3oRpVoQrmYhQGY+ickRO1vQi7tLmVpSNzrYiU8fZoKvTc
P9fnR8gKVc9CqUgLMqny9iplYifCR85/VUnnaq0hgfYuSrvBt2HlDiDZUaElOG6xCqKdv2FZxf2Q
kJyHRJfEMeJNBkJ/9b8pvL1zxqo3laletiUGKYzeh/vHt1ZlZhkcAj+tibWqaKg6UinG8ipyACW2
YHOWfrkx888xOAWOi5Fm19I4h2yK3x7cLI/zuCYc0UTyZjfwpQOro5ZUpZ4WIUmbdpH/SGfyHQ4d
dJV5x+pxqXC2DhVqK2r7Eh9M9wJWwxPRwodTmGh2yh9txtf8eXAMH9W/0vL65yVyy20hkTphWyqn
+Kc/VnpTaw4qxULcBNlkw2I3xx3dGIHurq19/wj0B1tdI7uLhnDk2P696bNk0fEi9zWYwvIPyymA
Wl2P8pMnf6M4O8c/jUs3bxCpheTFXjiUb2cxjqHEGbumL7T+t3Tyq8NRnNZ+MWXRhfRCFclZfd5+
RhIdan7JBNM0QSLu7LJdSadtsEcLPhQ6rMNKgkPpoPE1w40E3x5jiMxeEIw0vCVOxL8+HWRQWVl4
W6x9IATpEXZI5i/XtVbJnYWYwzGw8MrN3Vgt9DeVJ/HjKC9iMw+vFFj46akKIxdnnWtQ2ODO43v6
92TbChwRL1GL4vFlLDRy9WUKCg+f4ZW5iv+/rcIoGGOhSPN/H4q3+lXwUUsStkFGHz3R5a9A+qKK
5Ke+e0KSNK3a+4p9wZk/iu95+UKNeMPRn4SuUEsmcdcsjJYX36TGBjbOi7qHR/a4inIGj3KKahT8
sQyWvv2AQ9VwRpMzQv7uL6PMboiUAcDgbUc/rN0oLxpSbM68aTFxFy0LD5A2cXbJNRR9qAJCn29Y
bPbDJG+daKpeuWIxQDlRgengZWCky2hlAR/Dj6MoFCVFMacqrJHAjCup3dbsjZ+gMoazXShDpTOa
jkqO7bXPJ6lTSxy4l+kWy7etJorQCm3deFg9Am8sBoGlKJYunQAT9isteWKKJSrqJFXQBRbZmbIc
E2Hd/f+za+x1e7L+AzEx0mfMBZG8OJmIION9MDSd8BBlMY4ILuJNOvwLBrnQ6rpKoyLgoOid91+n
Ftqq44Bfw1jL1I8tM2EUwQDqEsbsA8dRqJ1oEcpG1F8YD9bd5qe0GJm9QNfdAmEefGsLJ2LlnR0R
iXRnPcmwgB2s7lkcfH6RBdBQnOIChTXDM+MkhljEjHjmmwqe9oXIih9vvPdjl9QHC/yQ8m5GSrM1
YrRnchYQdpDSL3g/id+t8uda/VZ5I9C9y/DeATStlDYmh0G4CQRkRD0/LTxIqhnkTN9EujoUoUoX
m6TW9PDwu22exF4jGHjvI6FYb139apULlusGDyULkofFYBHLid/MTzTC21ET8OKxfkx8DZ/rWpWH
exGy/RF/PqLFbMPKXZmcIv0oQZSczPBeNWWpoJmLBYyxvh5tviky/Ba19l31jHWFGAVl+i7YVkrj
ULAUMgHipLk37rCp0Edx4wyVYSQ2oCG+PdilYXdiH1q6U40HAP0DngHPL9UTYgz2ALbIB9caRsAz
B0WvzN5p6l0O+CAtoJycNaC8R0hanR2QJ+HVAc6ByOpjAPpTmCa5c2kw16XtecqeakEaxncMK4Or
KDgtO7GK6otnJ9P48Kl3Ct9s/orM8tCm87xVwMnsipJb0e2Jjbe5vhpruCQNEGalduwfbv3uS2rY
36yTvM9H7kH3gKhB7oaz/KT+WDXXXKR5TuHB2gUKrbL95ExIcO07dGG5KJW3ftdCjuCQoc8ddJzC
91PVtGdpEMiAX9Boicn/rzX8e1WCKLXMMCVxc2YmpcA+0nRnPKAJelXgRJM2C2uB0kuaFNvieDnQ
eURTDc0Q5Cl6PHnPkvaZXXusFVGljtUiqV1DBentxwRZttlgOOAvGpCExlm3HKJXEDFNCZLn3zdU
KQDJpJyszMBKvOvnev8GJk7OdKkEnj8NXb/Y5pD3UUaqxmtW0ce30wx2cwHGFU5UQYwWoiA2qx57
3lZFROotg3m49X6vBqhKVAoIyPISSoeHpufdKacLqgaGtrZBAkWXT/ZnAL15p0Rdj3C9YuRX0bEq
cFR56Tj6D3mpRm9WM6eZ1Fu5veGSiObeU+w2NSvQjkYA6RqrD81Cbd0YgtO9nDjLlvGsFCCVFbtb
KRiIT+oC0/YsVrSoKoubsa4zP1BtIxiAcvuv8Csong39k88NhRG+oy5FS4xMo7+EkqypKn5epx2e
5WI+yO3gp5buWeaBgS1VGz1CZewVdgqYGXRhHOXIr4mgVrrxtH6AOAGoimbwqOtuBuX2J6pWc3V3
MnYMEtSdswTe4uszvirHtNrZYUVCKaXsjsOGT4LFtNpjp3CJT0WRNdyAKFO3mVCDkTxfaPdD63Ho
F2HCTTBoTVNmYXo3hPkzhzTkqpI4HRQBDPXWpbjChCm9m7kGE9uEFnQZtWhp1McqnKKPK7jxVGbB
Sm+nLH5IzSrNdy0nGmV73qUr5aEKHMTn9v2Du6khg3Qxilcy+HjdyxX0cP1n0aN1H1w1ciYvp7bl
Yh04kH36Y35BtODTVQP1LCWWEZgaX6gfKzWNhzMdzTZX8ZpACHCoLbyaU2H7JphOVJEaHCDH23zX
DG2J/gP9kaC9KMVktRHBBf8XDZ6EVTwAcp4A2iknBp7CR1Am6hQPfPOUyjYUR4vHjMGCW+u+rhdv
S9N++Ej1UCFpff9arR6Uz7DK9Fk2ePIHprGKc0+Yn0yL/rZG1z0O/fY8yx2gxS6SIw5NaoIGV9sz
bBg/MAmte6bIU8Y1wQsJUxNJw/w0IHCgwbaeEmQ1hvRVQhWg6kJy60zMBbNTx4v99s10BdM0kN1W
6QXC8hSIuJDo2nZqb0ROazKeLsFJR/vygtFlIH2Y9nE0W43pVdlk2xHuCgEmCZ/nczDaqsiI8h4y
voRh9uGy7C/eofaT5gt4Zkwn+zrBTcYkHBQlUD0lNqdRV+HIs93mWw/l2sO4+4UQl9qv4phV5CH3
SbfGPhs+gdsaGRZgvXJyi/4pcSoiZ5/zdTWESZnWEhY/x2GrQOoiYx1aTkjZ1C1R1y2SrKElehNe
CgEeeX+0KUPcxE5fk5v4iwQoW3psYL8sW72os7FmB0QY3EQdl8pR0sM7dsKEt/tQOCOS5NBEz3V/
raw82FCgYlalkSeGwSiki1Yt29sm+36Jytp2pEmNWEWo1lGHIdID6wY1W9/6tKt0NVppXjq0AzFq
B8BgEPJuU6phsMGxB/3SCGO5GKj+33shW9uizW4LfB4ImH6++oUI1sKvUm8yqBIcv4iiCbDl9FWL
iwUpg7SbvrXK035XsLF9Uyo5CbkjHOLhGqV8dsoSLY8dSgtMwr5I+F//RmMNTyiANjtwvCa7+/Bm
ht9E+ZnX+1LeIeP+ZItxuXo9VlBMpm16vSu8LJoJhch7209g3Q5DsSqoLL1lU4uX0hoSduUrEfYm
g78xX7xLBo5JC2w6wb72hzOuxgRahTzoM9yPcY4MeoL0i5cr+F2eafv5m/ow8SEDZOHrnSttd5e9
gP9uSrGqKe3dm9/E+1jTjhitKC5kJ0rEjpRpZlRZYzi4Y37M84OE5zjiPnR9Ddi0vW3UZ8pwjJUe
XI9Tbq4f2RLjQNfZqQJJjYH+M8NpsMjNPW3+z53NfRocXWGrnLhUvX8bGpKLEccDnZy16hlOHsWQ
L7ZKnqlk5ZUmAYVFhCKutOMrGa9h/Yzzbd/JlaqdXHXnL9HLgemrAVjIUsYJRjmKy+wRFndE8cOH
WaeP8LNmwg8/ipg/mOnAyrwSvpde4v0OEJZnZItsxIK1aBdrMl/9vw/c2JLVVyxn5N2sXGLRwzfX
fqm5pPvpSkUmRoggZ0WANEE0Z6J1tiMlPGb2KVWuIFRc/8DCyXvtJ5ZtLe8lixJFTMUXSqYMgSNs
V9rEuaKvf7m+21UTWNZyhMXSwGv0QX1Y9/6JJ/+3r5u3cowf2SWyRVPSFXaPgmQgMeK975UjMlWs
wNCiTJLOE/fxWx2MjjahuylNsCqAAuhGFgz8t8v4E6ktZqs6FsIcNN7zRmS7HyfnB3KFPwGjISyW
LkHiDxae1ZSEhcj1pXtJ7IfCUV8NLk37sfgXR5uCQ9g9tMxn9mUYIhBV8wJp33J8IyeDn8fuLSSe
aGh46tSBO8GVfEINmuqyV9Y1Hzzp2EBjm2gM6hwjSWS7Wj5R7SGfsUOFzNO6HqSdkCDAkryZFhPn
/PJr/STbUL2CResWaXGxce0Oedtu/AHXZIGxdAWJ/mJMCljPQsp74JVq+HufCE55RFltEF7PpvrV
SWgk1yvermR7eUUpUcrEP3e1jrOxVI9GuN9NYSVRspmhGxoXGh17gTDLFJpqHGDXrTwvfawzrkLJ
bYbzu114+VRNeam1aLLsGOuVcQhN2JD+Y4A5ypnASznVGOpckiiNfg38h8D3hko1MBKUcmhGRkvu
KQhHZfBW6QwQb7eacvc1Ib+xtScA+L1F/brhcZVfWMYRKZQJHwGR27iEr/TS3iv7ZFZw+yf/u1bO
woptnkUXsuZpHROFJJte1WAvxJwXoi5zlXpY76/gtAdDhWDHarPG3X7DzunVxtcbzR4byF2RwOab
HxUQYxoii3+NkZA4Ay2jw2NiYJ16Hp/fLvIFf3OZcyakH3zFaPoPOZ7xlG4WIRoZK8FiLPLeq0+x
p2tEDSGgKxpgE6m9eOCebcCaycpxRsCG6WEw4szvjIeNE43sBlVYpEPrMvYw60O7o+TyBe5XhPe1
PqpfbLTtTxX+SFgq00CqW74uRepBoukpaJ1DlIay5iV/Lc53dW2cb7LTyTgpAnjDPaM0OyjUbIL8
TOOgUE+fjwgVI05fDViUDdtN4R3y0iLBFQ499eyWFPSVbdbqGmN/JaQHhLsYu4lMLef5udfQD03V
A4NoclMHNl0SFfsiy0PVb6vsJlMyUKiBDR2nhWV/QiGJ17Pl4vEj4BjKmM9l16j3L4QBDhRldpcq
cJgL9DJyQFG6mOLMTq7b8U+he5WWSuT7M2dBswuBrwuVTI0kmR1gunfDybCSpNXFftdqMhHkNo92
G9XU/gB+NeeJ8Cphz1/sj/0uAov04z1sogvpkoR/Jd7QfaK+X7vOX6ByL9SdcvM1/X/DRXAobhQ6
ZztFoxEYSf3e05/KSNiVVVFzhZeF9B7Tl+l6iVNhrbLgcz99til6Lue+JxggiNPT6QagFnU5qeLi
SPjQ7dNj55qEe3MkO+FxMrdOumPOOhnfP83iuIfRg13S2yJMvFoEFXrHULb0IVGlS+mXEcwPFG+w
sUIhHv7rYJ18KNNg1EIxwWIKsJJ3Bdd4yqpzxyKof4fRYWnsNDXRRwdbCtjh2cSITUfoXYV6KHFY
zcw5NRfsFuUy4V8nutu6np+o0jGGdRigA8omp2VukmcHL8v3fT5yN7Pkb2BfE2MvVvQ/LQcdkkzA
ZEtuhjTPE9FZnnkqnyearUnXMcUHzoZcxoiSLuzts6hqy4IM8GubpHKvrbOVzs8GH/qpF1OvSnyJ
cSFzZ/eMjbUtiXTP68VUAOnQBv+HqMyucf2BkH8I+cbZdy+MikJDLgTg/IgP6Tawk72Oy1p7mSOa
Z5VE4akaMQ/4ELbiXHbxHXTku7KwjMFzu/2WX0ys0KUlLyORV2QwPvFHtDux1uHIuBFWh4zhEQg/
SsJEHMkMHtwrDYPTnSDUAm+weuuImvp+UXmRxdRxnWtt9MRHwYu03ydZBP9140S5CivURDfC+AuQ
Qx7po26FcnhfFj+TTLmNqUWupLfILuqH7DRVTGXcWVw8Jjw2VL5RCezoMxbjwWTmHrHVGiNieUlI
3LgWI+nIRglV2OPtPuVceG9M5whw5UmEFWTaWNjl5bygzMbEUJEeiMj/HUlh4RtMxvo3EVAMxbSU
aK11ALBPyg2smUZ+d08O3cyza1QeIo/kAcAK5MFHotUQ/sk90ZTQE6l7AMmLJ9b3OUPxvjqpb6vk
y7MmInev1JNhXAhXwqaEia/hyZoV3OLp+boz0a3qG49mRgp0/dRfZDCEYRYwxMs9U6dPSQw/Hsae
Ji7ydG/SyYodCJ8Oql4OVnK8v3ZrcC+MGwUiU2jfhuvlkGLPaPDDq5ZsAEGbzf7LZYhb2bnHgnut
jD69OnoIzI96pMc9H55kTYPaOXBQ52RHCw+HUn4lIewbXpdzGy4ljLC+TWnRyQmMj5+ydX479Evs
HML0w1vkmEHEKX9p1VMxRgyxA1ov9v4vh+NjuPUV7J+MfiX8lbIFVOV9HUxALFVYyajjdUrW4fUD
4ODpWH8zcLWrzIKVgkW03I+ZulxUDehCe8EEGgW6XEcVIMI6MYqzktTs2QtfDvDAmWVpPEGBsoVb
6VxGBGbjiwzHPVSec1aejwSChp2Qq6XCnR7rKYn5OIhFHE7Astn5mJRXrFLZ5Vc8ANImoRtkzmeq
KerIyJ8fN+VpXdx/0dXLCQ/HWNyCOTRsmIBkVFVUHW25YQIkw9h0MLu+RvQq4II1Zj9M6YElyJZl
OaaGX/bNHwReRrpiuIOslmn18rXRCqGUEPiiLwPr9tXi0j7Hgu0ZIenVsnuaJTXFO/JsO4031D4w
vqwAt5+lOdVmidhQISSt2D1D8a5JIcPxt7q3/pezWPzlZ/l233r+Mlu3f20CY3yC6Kx5tASng0v0
nZVRmpxMbE7ljGTW4xN+6WA7SormSvHyPkwtqmyRo19FlKdD3ZdfLInno+ZC/3lT0B0iGyPI7DVs
F5DYBX2gBeiH8trUwaFlCg+vnZ/zlBf8Bgxh+/KVS4xkTw6AgZXHYg2S83JxK+Sjj+C3KT99pkxB
PxBFEZOFBuqRWAaAd4yABz/VuBjvRh7Ss3lOze9ENHCOL3KgZmH/9TV1Yz3JlFgLFUD6yvrfMEVQ
UlGQ2R22GLRNOIc4179Riujmcf5/nyunEOu1BNaMCROpnH4p66/IAqy3VWT7zMPwUYixmS1Dy3eo
YgYXJc20p0Zyfb1wyguFWKNgvTNJTBJNjlxv+QBx42eUwnRlNEC/rXRwA9uv57NK1SklvlWtJhUE
sRjyHK+IUFEh28i1tRfnyGZR2i37vPXUuk2JDCfNSW3vJtl5QW+UYLRmhkO+LIYT/I/PPk+KMEWJ
rJnf4nCH7EmT+zB50zqKAFSc+WxPzB1+SyLMGWcJxWkERjPhEK3rqyt8HkHZsflBkRlAlPPUuQWm
vg1IcU3YatDN+8EpjVrK4QqGkMYNiJ+giJ66Hf/6dkeaed8pOyx8aOYWLz1VS3d6btqCD8nif+IH
uaYgb60DxYBjdGEyD4hDgFxdf9nn2/1TTB355UY/4aQ1WK69dSI5wpM9TAsZqBwQZHCGQ6FuITbN
fnTZNvc79lDUlNlxKf3WvqoHd+L8e5WVUkx5TMXC3zBf+JLltuDX73htIlDcxzPotivOBDosLdvA
KiIAJr+KEL3XgrD70Yfhj0MYWHpGReTtwTVnFRXDY+4BClnHi21PJJzNVkGBsQahJ1kMz/rzxH+c
pgbL9q4wQVqKJn2d6lr9OJqaimJQSJ7EOuWRoZuwMMSARiQWmO+JD+JPCuTX1X/8tlBtlVtu2YAC
jvSLsI2B/I56wLstKRIufB0p+RlQq0pyiV/PTzypHuc8Zqe1TiJA2JfvDUDuP2EL4U1Cc7xdJ0/k
cbkBRiKFeAtoyfcLKQroUWX/oYJIgQt+V1SgQsb5IAn/NHwEd4WvorqjpE5d6CR2eIl5uDnHcrOK
pUYTZDx6rV7qaaaFMXLiHVoLEBfoAfcQZUJiJbBsc8ezaMDOLvt2wNhSn8cWIY/9Dr/k5SGxMJxM
ZtI4UP5MvxhKoJc9JucsxjtgoQagxneFDIXbgHi7wfuVFoVFfEIjsU/U6777xpp1dgS0LDn7wOMM
uT6d4k+J7rU2Q5pdxOakJfH0o+b1FANthY2y8b30rwQHhp/Fuq+ohn7GDu4E60keXJz2VF0S+coa
HMU0ca0IC9mS87Tm1c9hNBdxDa8F2+JkUe5+FubsRYIoWLlQgnLWcfhFFgagWHdedPs3A+mkAIkz
XHuION4vHnI2SIlpn6TJzFr3PzSXVLEnPqPUUd/x68H0hXvD1UDmjamhTqRgaJuoy8BwkJNXMAxS
614qpRSY0GM236EX1UjE+Zn5SA+djvLJpZfC6VY32sRgOkSSJ2MyAJC+gfCu2T5TjCfgwcmGS3UK
LjI3c3Tr49LPt91HdjykPjbAecYFLHCaL+Ypr51o8Y9vVgV6z8pIRnB5Okyj7J1AVIgtFQMFz4i/
6ffB0QHuBvqFI5FIDR6ka5W3Dl+6066w6OplrB9mki2+82ssjhJT9HiglZhn4sRUIEbBfNH5eZ3w
vPMRalXJK4q4h9hAxEsJHPA/6WxXpSRYaktrOz53pWW0mTI6E+AmA7dfb6tKdtJf7Wah0ehrFuo7
k6m1ZSs1DQ1wIL9xkT3IMtiXt3+oWVipQlYRM5HhPC8VR2hFGmEhtrBQ78y2ZcPoqgCFy50D3x83
14+pnIqwst7IbCSCzkn+TtGI5Li35lwNSQKZT//t6o07+VfYS7SCJ+voDcBEdUW1aue2dD9efUvt
ET89OhMLM9GYwI9Ir83wpQ6WJDWwLz+ZTJmv2M35Yb+/XHhaK2o/TrRmRXiMMBXFViuNKzuFuF0r
AUy/EHH7pR+eerITZhN1x/K8QjA6wpfAqGzBnRhHXiHNnCvshIQKCORaaXg2c/MvqVJmvoeJvFm8
rn9+4Z/dkpn618gdZWWkIrEBgC93Ji0rWDmCnTyXwTrkTNad/H4lFeeVj83AE1ClX7SR/iYI60wm
+yC/WwcGmwb2bK2ThMtxOYnpKF5N0i1RkaCWUQyRR9LsyOOfFFKnARpy0RJaKGBg8JgCaF/+V6KT
Y0o+P9KgvSlNzDlU+czWAOtu05pi4tjyia7VaM2PpZYXf+VA7afs/MLt5ZqO4gfFGc1o6QvnHXZZ
vZ4dnQ2JNsk10110g9zBAajD/Hy05Il/dqLjgrvVMkO8lZYrUbWEhrkls6I3AjHwEnbe3lkXzS6q
qOr5einpZ47PijHqsKvWP+yE3viw6rLAgB3XnPhgL3g+WldEKcWeRezQYb7jA17rBUb1P9cua7kH
dgMLCwX4UnrkZOsG43H6exHAd2h/vGyzLTrUnyvDH0HQp+193ihAABXYE8PvPXfcpTg1RF+qe/xb
1VjcodETiCoWxGWgWq4d1f3Y/zmouMvdmfxDyMQmkWfuNqOxzhLhexVZwEtzUOjpC1pp9G9Naq6v
yMHbf7alzFNjcqGrrkdu/hMw6sYgnBrzpr7/Ju/DvHSIC8vtdw7NJOYFSyp/Ti1Z/fNa4hDp5+it
pzxfCInuJ0zq0F2XHLac3KEZ+9a7qJSM3xQALg2oM+ztWfWyUyzXqlMWd2eiJoU3uMOVQo5E3/GI
hU3FW4uxCshBTgfLKx56CWU+CZcHze5kZM7S8lb9DIAdCmNoqwlE/lpWiQsHIK4KDD8i6kQKwKSn
oH+fDBdh7gWepCSWG+wJG/TmCE7aUXFINUU+JI6rffvyJgaUXKBl43JaPvNsmiTni9TUs+JuOTwF
+jmJhC0aA3BFV0yh0/+e3SuAhNzxv+dsQZ4HLVNRjB4LJyOFhm2hO2xA/9WUybHo2CKGuT/pKZGr
wVNzj86EYSIq+3eizO92m8AKKhVXbwpVvC0umnyjuaDbrym17xX1WTqtMszue0eHyn28EBNfmN0v
Kpq+WHW8b3McP6pfPhE5lBe8xbZqgy4mET0dj1SfabGXtFTecsAC8wUb7NmmPQOi6vi8zhpghqv8
/AxumAD0E5R3TSgOZBGZDyTsAPeh15j5oyth6nbRYYLj9rM2rRxuU1V4m8iS4Bwpc6xwPO63t5Cj
DoDCTQfUKokwG2bVANLKi8AJOX6wMj3EdjfLwz4e7zSPPGQuctW/ubNVN119eFbl14eQtAox7pPO
FC4s6ctrCUozvsvgfuRIC33f46Qk0bRgxFzHG7qrQOOKQ/tYW1TQfbN/sn9bD4A/WwzeeHOn589C
9p6yUgKNa2sn0bGCF0dkEwIpuFQUhK+J6Yc3mb53HjCPwiCNNXKos4vwI/W6d9h2SM+1LfFwhbBd
sgpXa+ArkMrdT+nGrCmL1E5MvIWQjad8OPLp2C9gXFa1huaaNquw5kfVtfS8pPqserbL6eOwy6l4
Kq4zjq9mIQ4WvnFERMKh8RBoY4f4MDyY88LaE5OoTSXPgrq+WeLinKUVFZlzz65BBMUsGcKFVCt+
udhkm/NkLgYjg/VMneOWJw6tjQECymW6BfQhT4fX9FtHtEZlzpK8BV41ICv0GiA/DIdTSy6n562C
wCZISvkCvu0J+umlXPPmwSXdQHO1hFxCe2qSDrfea4Bc4wysYzFzDhwDxgTk6pVpx9PD2bt3AwqG
PQVyM7LRHOfy+VA0oXk1pgQwwdGveiCFl7sGXMUFWxabDwpjA0Ku9GNu1QCt9DIjRsTereQiBA+1
mZyxAxDjBmWA3JK1fS7qSz9W4pc+2GpmoTs/C2xb8oomwFwo1Jy/OEpn1c6GN3LSj0zTXh+uAINR
XAa4yRrLF8brs1HqDUM0kl7d23jVF1Ym6wWmuKeuXFwrsmom51w2dbbWKffvcWrxi62K/Xec1ueK
vukgI6hxL5K/LilJYvFvHpQd2GjG5X+DjshBHzV4cPFifRIbc3fI4gl4bw+MTgD8k1PtphFRzHOK
G1QhNiBWhWBexT+h6SQfiB0bdvQvzoSoYhSKaFWmANv9Vhk2ZcXfVNs6g3quM4zymDYtBTLv58IZ
ea17fb1MJkkgZ9d1UQZxa7WQbGpGV8nVrrEiX6JgDZohgjyyL+IJpSnH0BBLVrMEeYRw2hmQAnpP
bJsuZppSCtQBAAaY9yn5Ei6pOkkFvGDXQ6Se79pcLq44nZQjpjZQ0217bCsZ5isgPtHM6A9yUV4p
1hjzlOvsFsRg0ZdoXtNT8y+JnwELzw6QHYfKbM4HT+TkZgyYKbQ4DdEJnmWbxPcjw5stdpbtek9j
Voc4JIdLT9YBsrmgLFpol1vB3RyGnd7dKFTaJ7CUQMXih4QCFkW8rCHjYSLF8WOF1MsnFDx1QJK5
HMZvAS0ivp6IOOkwl9VRGH5bqoaxlA/VyU9JREw3RWWxGswGv4hU0HtfUtwAXX2sDX4IsATjeZMm
JzFTXJOPqGUDjNb71evoXFHU+HIJDRSwHk8N9g02N9TxlI8bc2sB18k0l9tDHOmdizKBtbZTjK46
V9a2OeR8bP+ATsvw2726v+U7pV3KMlXk1KdKdc9QWnRXKA8i/3w2+FN1f6Adozd5qLIgMK7tscD2
B2KiBD/2tXU04RcWt7fd+FAVTgN9+WJjzxUJmFpECMJLZOWcNcfYecFhySifmPNxszLFlX0MIXdh
xohrTyTXx/h+byjQkN3V465QnkM8Arfugj2RWMoX7xitbgnEbmVqfdlmmhKodabFa+vN27COxBVe
82nFIF6tBIfCa8aOWQVH57Z9Ah1LLEOsB2VkdJT41of+41TcYlMUFmSHsFMl4SwB8myIGhLZLo+U
Smi0xhhIlCGBMImVxPJLLCJMHLwIpcjeJUOuW6XxbknA2YJX1MMTOOlOCkBZ+Sdbo3/UUHdhqKeX
Q2YwIkg7Ay+0xZoBeVf6Q0UqcqUslRdbXPE1O9bUsxMWjyltVtxL/bjkkamAGw+DyWWKD9RpisK9
AtEV0Z+T/p2uolJ0yuJnplRnhGKDtzFOE9k1PUTVDmXN1HJFD3VUUnAo191TkIL/SK5/dki2cHUk
mFm0vwCOEHpwV7NZ2Yj8Cp3sge2BQbIO73PZcZ90amUJXCzZQtpZstsdUGKwYrJn/PA4OKGqoP+l
FaK4tDo4cxJdTz2MDFAItE1eBTSdK5X5ifnkUJLqKXHv3FyGVe0UIRQc0iJc9svW/xuaifGry2fP
HzzMGGCT+ktDkveeTguGGcD6+rYSi0NgW9MgFyteuoaiaDz944HltjdPHSDCaDjrmv/TQpbtEPoS
VK4VCbAyLGK63R4vS8/mCYIkwYsKInLxmcDqWfS/dBy5/kL6cC8Z6SgBVAxqr/0rc4xUnA8qfRkZ
tL77yvtKBHcs+cVZEi/v58T5ghHf2dVZ3Bridpm/F3S/RWt2iofWJ+5NORNpgU9LoslQcNxsHUWP
72LGGxOo9YyVoLnhiwLN2GNyV9tfKyaVkjj1bxF8YHbVadHuJ+G4j7/lCe7EJnOJx8g5K+WBgdzQ
xjZHCT/eh7N5BYplUUg9EhNIz+i+9AhOMlnCXt2GYwKOF+SARvvMlFqXjA8o6iYDPLwyc6ysTRxO
ZdZ0yUHjkk/4hhWBsticYFjAQYkB69KmzCQ8IgQ1pi1h3UoXXW6Qr88ngkyc+bjVICYuxFqvlix4
qS9HMng3MRVqyIVcAwXbhU95krjUdw92SX98U6b0q1TE5wcLKzJVm7o8pgZXRe2p7WyVsZQNS9lg
dj/sz04nsSWRUMN8lR2lNVjrD9p0tP5bITia4h7zlxim+A5XMVEyocZbX4Ff37N/8EpP75mAEEw6
38rJ2rysU17B4//yJusQ8LLjyOIjs9sKTqEnKZa63InjUBSdC3NpC+5DFv7eygSaMqv2Io3TYSFX
WgVqe2mQw0PWS3gyzEMl0S7YUfSwPcoi+x8ks8xzrBEviZkN5qr9kPPShEI9Nty2Icqr51CdeFR5
kiX5Pgid/C/kZpJohUy+uiq4QaGN5+i6jA0U9pc2gfaMpLlQwkm7LDXeKKPmVwmeRDUuoX053MXY
QIm35G7phAJRfxsTYRe1MuqkZJ2IihQrpUd7WWS28QeU/kedz/e7au0aD5HEArtyoVUp7a+SCgck
d+8/9L8etzWSMlxPz1AiJrGbJMHAU10cfjT0BlvwvD+9uhDi3m1OTdUwLLVeNLxG+VBg+Kd33dF0
w5AUn3Jn+TvdzScZTWsYcGJY9oeIRyH/FSir3A2IyBQs9AZrr9NkQezV299gdTRO7k9CILYGxDNp
1oUncOezieIV61hgXD9Dw3Elb9Pg4/VMii/amrrw+U8DKIAQN4+b1Z6O5XtTJEHeuJIe3rwRL5qA
ADkBEromRF8+4OgMlTIynLvgCeJwCm6vLglSZswvahsVaZxRghbyZ54g9PhJuMfIvu4WM81whVIQ
QClgulH+SHqvoAKbu5PPHA4VTHst8iSYmX+fwV8Qx1k7i9wjFT2uTwaYMgiXbZY9m8a7G0rFKLku
yy5yn7RfoRLXeJo83L8oiwKS0PSiuGUp56utUlPRvrxazuGRU/1cN19GFV5dTE/v4m/G3jevSB96
VZ9DDXMC/7u/PrBHn7uD+6OFRR61wDhKu8KGUX1pVDwvyGYzKMEv2DTeGzeB1GtBp6GZK+eRCwwU
u3k1fzl+mbaa2TbALLPwq7pM8GPNsof5g/N7HCdIKOMWNMZfcZ8/wIH7WXTJawrW5JUYYE33beig
XCwoTabqvqJd/Efl1lZOxp6goYb5S/aOCMCJnTpqa7WKjRCAvU3YPKNm7l/ybHnIfS593fSWw/BE
npPcqJMPI6biOJV0B03fi8Cb0xHWogaA8uCoP//Evtts9ACBSAHkjle5U7Tjq2DOdCpPTbftDNLm
zOZxGyKE+/PfEeiXYJQzhPpwGlBji83mGzMAEpxJrRorKlRAqYXF+qJCsjCb2NGWpqpjDdsF5ucr
anRi1yoCPzcc+vFtfZuLOpKX47delu6KaIKVhq7kULVtGpELbGofqxs8aVvk4ZAF3Npp5GHM7M3d
V98hOEqMilDTNCeZ4dvPbWbTPfoGyqHfNs5QmPj7CAoHKhduUacUO+nznl44L9XQIpo+kB/TyYX2
wurwK8owX053IKqP8dm0AUC2ANQ2I71taODZY2judCeaE5+YEZzxPsyYsFbc2WJ+/uWXcHFX5s9W
KklJjDXNrC4rmRZchu5orujwBYI0mmF6yDClS4kx9552OrXHBkgRc/2SzkrIS7hN1/YuYeYspm+A
VH1G/pQbnSf5PunL7lafWkpdpupsTH6dWPM1sMpczLz6Mph70zWFus6qv2qYLGXOqbQzADy2KMlt
ARIRktiQQDNdr73iUmkPPdcXz5YFfYiXt60qFsIFKTYSjjA3mKxf1v2TQjh7nQhvogYAyheAPR/Y
U+H2mOK9pfdCnSo0gN70dZtyrONBbWM/edYdMgzaNud0CWHGcC0JAgIYnqEOxDOsWzTe7K5IG0Wk
WaQ+tmOBpf0k9IgLE2zZV2D1QzsHA9Uo6U9KniA/OBY9VWdqXnXDe2jqp+dlYvUpCmJBIOL+d6+0
oLjiZyktlAkUw2Bma1HX3kyfDSwrs+bivOeOal67ZamsdQ61E9cbkPiunYKWrfZ9P6r3iOAOGMe6
2MwJzkgtk7nXNRFAMIlsXXI0JEeTC+nViRg13j4xzyHiJtM7aK99rNANkZ+9MMySwqANG5HAlWQh
sAZPmAg0m9Asiu4hjds0QDBFH5zbp0mVUJnl8PLX6kFDveQTqAT5yVGeuONzonr0CVYJQFL1KiI+
pKLXYWIns4RFAeI60Cxv8MRgkwRQlLdsC69QsNIxrJgQn4IQBr7B3aM4yxhDfwXJAxWLNrJH80/X
jwvfyVuwPEMgYtwcBA3VCFw9ZYS4+JR0lE5jtWPCT34NiX41oxsUR34NnS4QwhSLMaBHP1P6rLq9
ZWogwitdKX90IgAVGJjA9fQBXo5a/g+XveG+F331RIKo8EPPpEOeYPxxcjbHGKo4SjrLviDLqKCB
AvH2OAsOcTtRLJ9Gv5rDShPnbuWx6PhyPo/8yHgPK9sPy9qg5yqFckO+XGhvaW5dzv9y2nn8eCv/
wCt8DZWrx5YasEV84ErIek90cnpFfMnk1gcDfakavqS5iRGbrvuqEyhN7pNLE24P1tVnj3AggTEZ
iTqB2s8LhTihUzVae2UJZbkIdfw1dJsQa4DZGiKtPyClYWSGPlj+KmThD2QWZKbI9DFQ96eN8tcs
VZ79pkAb9M0KY/YdllZ8O0xTNDr3w+CsT1iCMvFmR6g3ZX6Hb6CHAlxfw+EVgxsvhpsd1eQweT91
60fcUy/DhO73hYfpIZh0R9beN4yfak2/es0r0mAMLU1yKn3bPaQcV8EgwVN9cypwAZwfBl1B12fK
rZizuiqdc92L3S1sLjFoN1wtq/R6pHterxwiBvS+06Xe/CqfvucYzt0OTXHipa+nqmRYYLdTRlJk
GA40aLO9SbV4OxXFB7gl0H6KUNxSj83hc/+nl2AmEXqSiyu8xMa1NU0g/Fq0SyHk2AlmnLybiXY1
fWAW18nourouolBUzANb/a0T4blPc98V0ZK04QTURXW+RqGHNetXUT1uJEyeGQxsgAH+HrqJq+FF
epT6XaGrn7SBGwnwkZMJ6XwTXCcMXIgwuQyeuVhiEM1rlXmvnNxm9Z4oZtpXCjXxTUuwmvBUmBW4
KDcVJ/curloD6LJjonzuBP3cQg+qnJvihiA8/NGGcsmadBP7TiBELnSXwLDzsvtuu9OLqHc8o0CN
BpUta3gz/2l0LVrGrQ6dz93htIk7b/3BKr/V9/z9vjvGa5zOyH1mnXerEhJJDAa1wB3/+HIE5p1G
4vBJPOdJU0nSCoS63fdquR3Dbg8SWzDSiYJCO1A/Rap/sqLTFvTi1JfKkw/15IeCBB36Ueg5pmns
9UKsNJ/ALYonBUAQv6YrLCadNU3hgTRHoAA3JT/RF9NFJGjUhuzoTNOwHRinvuqAroWMFiEbwqlW
K7dCyonL7faTaHN3UYmgERsRtHaBHshdYWiMER/uOiCK3uBoq1iXWDhXKVFuwU50loG2brUgX8w8
+5XlQQv+mM380fnuOzXp8Na3pyCOXjZbmC194wdXH9WLBq2gnaCObVlSuPY9WYlLcijsEGed/Uwr
A9fDXQewgT5SXi7HXxrWlXhCrdU+SHZ0RUP6TTZlEbAzF2qKweE0ErXz5JIpDsu2fHxtAGiKE9QW
G8+KIzpgpNZl6PtmuJCKTIpM+K2gY4/4YTozzVn2B9Kv0QqM13Ag8e/9Jsn4S4R2LKayNh9ctWeE
nYzuw0iqRv6ZkM4rnlEYaAZzmS0+JzYVGdvaFBDKxs7grARXARDf/OkmSHCa9pMhwaSyJOQbda0n
gtPYej2OTXbMhu2/ayJOj0WTN4o5LcRH7//YHhottlxDrQKNhQ/fPnsofaU8Yc4wEgByz8TVoxSN
rZ4S+gKZaPEMWjszqo31sQsjjM5KVhj0A4A/q/OEMtEG5u5+/wFJQaBfN4kTSsaqTaKeA72R6xzZ
MyhB5FsRhdM+du1q+q7FtZ+rAytcGxITZGNFMNnPjekgQmAwz0G03QtewIeAtJvk9jYiCW/lbVYb
j8TLRUpvszgG+n3fI9WK3vTm0Bxf3fW2wJT8GpIjtbfVoEGRM37UcTaeZ6OzVwFLXBBJwm2bGGfE
cSlSu6tbhp9FxXF6Bh1mudMn2KfTYQ/6SKl2mhoowN6Tyse7izTPjHSud5oUFddesYEyC/yjKBeI
3P3soOTZekw0UpoQ3p2VImDJ3nhWGOOQqIui/OFhVEpo1/Y/J8kPWISh/lhKJ8kbhI28GpWB8nmt
Gs0eYPjmuJWNm40HJq8993DawdaSWSpGyGOqZVSQFkol38PGz4nizAdBCcbxwDug4Ao1M4nuTgXa
WQw53k2KIHDXsOw+J4RkjAwkcbqB/lf/n8hkJ6cB7ZoZT6ov7HtqykaREt6iKS8CfQ5b+IEoWjZe
64r4RNz5C3ow2J4dKOylu0EDl0vBryIkkq3kNCTFR3qMAFilKA5QTw3kHzkQEWg+XjJ84SCS/qYJ
ka9W8UK6Cq5MAGSL8x6TtoiURMqzZIOfJZ963WF53ToR0TF8cY2nV+Hxati4qOHFo03BB4UsUxrg
ZCuMk9CJRxsU7k1+41uDraj773Zf9/Ej2aKSPRQGysfNYWhQUeNv8oLpBejEsznytyjORhW2KTN3
Bez+ziDM2t02WrSKfyJA2E/02yzEkN5yfcb2xiAt5eJ6I8QbNZ1iIc6BDw4Os8W0nrjdQccp+quU
Iqd7T03OPqXflL9Ds1PQLOA4lNHr/Wo5WX72GE4dF46G7AOrJfHKvQ5mYPu5gs6hkuTEw9KGBgnl
LxMXpp4LqTAxguNw7j43NyA0lN7O88AtQAnrGNMczVNJeHk2eHgHKschmsCWeCOWDLCfuEwvcJsY
yL3vatmda6RolmWtRLeqAGtflABV9sm65Ese5f+Ht7LhXt01uTzlLMw1cAsiLQwnS2tUOFDYp5Xo
XgphD5IjfnsVLF4bbOhOzkebZcRrl8dbbuCgkywTWgXjfZe0KR703Ve7Btqbay4tvqqRN4StsZvb
nwU8Gz1JwkdLvj6TPZr6PFuiSD+uVOcQgH+CIueiA1D6fxeMPtn/aOnyGkk6RIZOT157GA7N/B6D
wMbWyUt9jamcWUQUNGT+Fu2zAD9vCJBbTZEOEkMHnvUYuhp5A/sGJ4OPQ/t6buuf6v0oSMPQ/kpF
24SjrwZkeWFQ0Po+a24QIsfCJ9p4nLvVj7oC8HxqdS/ufWXA3xrYheE6aFn1zkFESJJYJuk8V6U2
LA3btiKt50FbTnDJfjDE89Lrc1MCVpkeCAZuP9Aghc78zc/xdfYP7D3VAttSJJ2jyE3kflyPcarW
jtq4YXLc9h0cTQcx3Acr3M4rks/hJqRQnAYMlsfMJwBhL8+qV1sMEC54jsExPZdXRD5c1Rqxy5iK
CTLyJtWYcLB0iSrhQ+5gXGSIEJMg3eUXv0PRfgA5SaS1MZLvFFm9nKZRGwKG11r5xSYcUhpoxpwX
JkCL1nyIi4E7amfw6C/MX5GWC4y1/OkTxargA2B4rTnjdSh5sLbJ2X2v5H9z014/vTsJdHICLdTF
aTTSkLMSS5hy0wgI77YO/1390pGjLKhDh2zLI32hIaGeNeB8B41R8xsI3wkX5UxxOjKcYn7Y24gR
Xhw1VZrT8Qg7u/xAPO0+Pb30F6fjcEb9JXS2L4Fk4pzJxkxs4cMk+yc94q4ERLV0k9YPpd07HnL3
TeAII7PQB9wl6GrnDlxHgPeuqFmCl51bWaFhLOOooUtVd8s7Af54evqdgtYLanbQ/CdwWVPvfx1d
JZYClz4O/F1ElXZBhKYlmtkE8Hvbjb4rtNX5ZHwxOLXjqjYPK6kl+ktgPJtmvd7ad8HRVpxooabp
80i6Fb514vpoAUh+HdLwbS3Akdi73wcp5zEg9Zbe4nlyjZq0Uaw/GjFQsI7UP5Y7+JT7DMpcb2F2
Ft/gfJW60jo6g6CDdTZje3sqyc1X/u7/IMgiWVIGrUdN94Eu/9qJwOZGjsXjwMvsuuWGi/D4LZy5
sCrOx1fpDgosdvC6YvIaxYN+G9QAO1J5qWYouy2smxaG9F1ulVGXNt0Jc4cUDuNq2h11SzT/QWPm
FDvHWFOb42xVDSlGOrqacLpe75vUzApDtrEt+5RPiDhGcExl/6/AtxwvMZDATwpLt393Uhrkr677
s3AGDilJhg1Bi1lUJruPKQOSmh6HHyiQYWmI7wgwg6ez2Jn2zj3HXnlzZMlRQYsFwnMMSl9EKaBw
vN3ZSpqX9Iln2v85DcRebCqoeaexL+zFfgfm4pTdOGcwHOfbwHEY2E49CtmOL0sugjvZ4eemOvur
/ftlaJsyjuaRtvGDHaX5N5gOpqm1vN69tCiNzUPtsi4fchx9fxqJmEvaovOArgB1o21G+FC73Dnu
yUVtn8QNTXC+jIy2qHozAX1biFkbHkUZr2IWJ+ka2t/F6gKe74ekuSw2zmYMGekysAJo1GZR8uaf
vpaNDmWKWktKLITmvCR346kr9/mgRUeCSAZzMObgfy/UyCLO0LV3L97lUFdaEVV9TXqLpJ9Hx52Z
c8s5XQ645dgdB865kCebu3Kd9pH2Ozr9ShY/Libb6odsU4lOXx4gB1ZOMRuXP5wDygudow/UDJgR
VjSJG3hSbRdqTXe+B6Mlhz5u7Nz+xl2Cd9A5ZcC6DXc0XeIeQB/+/3F73If6uGOdyUNVKYWHRCj3
6v6ssr5h0Ac2Jlo4JyqgRc2hMVL9IVmlXgqPcGngLouQ452ROFMkFZY21vOhtge3B+Y5l7ycTO6R
ta1A11xGZ3XyK5fwJa5I+kjM+9yq9/Vdnfa8pYGIeyIOZKNwcK6lsUFfQV+guvhczWJGMXslN/sH
6bSLnE8wE/P+Khfg4MtRoxi3XKpf9fAO4jBgvzf42S9s1Dh2r/O1CrkFGw1/Cbz4OMvsUYLcztEl
A2wisGRf499Kzdvg9Mo340CdmGiQmc4xi/y4wL0MrAi7WR+nCvkT4GXYXMKueY4jnBiAxzxhin8P
Nc58txdwRWPhjfjznZKLPZjZd+kKrZzcMJBw4VcHRjOWCUdCON4JRSGjPxxKrOp680KHI1xzFb1Y
hVTrznJ6bNYKn37yR1zPhx+ohI8GyTPoRH+cviWf+2nUqR0vzGcvtcf/G24nND7ybzbsvpPFxREg
uPx/16+MrOCgDdPi4zhQLGYWVo6AvoPDBQPMvAU3rWmEl9LrStFQRRQ0RQ2J81LNSnrCluy3x0yu
+Ar3xqutA5y2guC0UZK0z4IzjUs46WuGC4h8eqSRrM3DjjqlZGRZSSd07ABG8fxiPnPKIxezb7sg
p1fSyaHK7vFFtIvLVdod/TvwAy52NqPQI8x0MO5MNw5wdXjTvL+MElJZj99p48twCMXfLB3NVNMr
T5wbQhZSNE+4ZHQXaW1miJgizLmK9KHEmE2XypYSx5sP9907cs2cjx8oFhAFxYikV2kJuMyTQavX
is+JSXcHCM2/hVP1JVrc4YtG3Mjq1/6qheCpUfKqDJQYaseZO5NVQdIiaKVVXyD43x9rfJyjaF9Y
L5EDFXPb45MSFYCB1l/E6nAFLmnkM3n4W5CMYXsAn8cwksomuZRVeGohROTpU0spvaEpIG3I52we
SHWhyR76Eeioji7XpevH+C9Lo9eSZMo6KKLzuwZpbqg0rNiY0WrDLuzUx7UjA/NHCCZhed7E0l7Y
FpumkmweQm8FDO9jsEy3S0f3uiMIJtXqA0EYe0u0TS6/7X40/Te7tRD6Pgiky8t3RT1y/r4FruPu
+xQFYvlqqZTlIm6fHhJgYnTASJRGep0gOsVfzjzzpF5NlChfjyM+lt7g0xHnwh/6v9LuESGUodX8
qaghH5WWhSepXrVVZhxkDDfmhbHrqkg9URL7OwMDfURpUtdQXme135EGU6H59wY8Krua8KngAwVj
Ophr9WFh0Kpbs+e9Ht4rGg3ajvzU96hdbbgY+QzaHc3vN34G8G7kGbgmPx0BllLk/vnJX77ZgGNe
w5g3vs+ytH9qe/8PJ3kyU0ICabkKIhBNi9iij5hDose67K8CF/EG0DFo8GKobUAibpeUTrBzikb5
0Dq/8e5cZXhwv/CDiEIwShpkhVg7Ta3iWtcwCycGUFX98DW/tKCCKXjVgG/DrwLaJ/gxI/Sydv4K
d+PH/rAI7qoSwgvRL4R13qqsNXECVxynJADoG4smgCRhAH08xsABa9/gQUpX+1PE1snpHBVHehnp
C7DVj7OLg0RadBz0Bk/9Jfb4oNwfJvnMvO2vS67Qsa4cu2wDKJPH5IAQ+9bz/flfou5Zi9w2tLc/
d6fw7SxmEyDKd+Xne/rsmeuB3nQ45DWrQ7AStEbm4L31GOPZDY687mc+d/JGe7vESj3u87IGBUu4
oMPL3r8FYrJ+stGAiJQHhPt+mzIQYduHYS/AZWcZeTiBGGKanGk4C22A+kmua4FIyvnoTfOWC5Wg
tiGCYMtv346dZrYvXH0ZlohCTR8fmC7EZHZZsQ16yQKKS7ZNzfeu9MMJy7NMeKqb3g1rRZOWcHFn
xCuvdUgUwaNE0oFzTjNATHDFcQQBvPIyskOX5DtDopc0KkG74YxAXhOH8U7TiFqtKM/WCgfbXOyK
H4ILtbtAWgtR7zTTWWx10+NTe961Ug3rbOBTf17o4HK7HWBn70OnYRGy3avAvfs74KPvDIx6I3yt
9YB5P17rc9Ojz5h0fUzOObzdursQ68zIQ7j1+KASRZnkgBZZR71exdrVB+jiaJfLU8UNdIfxRS3a
vsaHHfpEx7qvMmnYXPPI+hXxqgoN4t3RnD+qyPbfB6OKIxxQK/bS6UrYfGiEdlffo49BEUknhwhd
maoLk4Plw3MCs4qC6cektFyfCQ2ME7t8ppSeqKs36QIJqJJ+6yL/8Tr9lF9BPjLmntm4hQPwmMTt
jg1ySMxHhx9jIOTt5Z7F/VCbeM8Apw9UK6P5mG5MtefsDQnOVtDCdA4irykFGksskE/KkhK12mHM
5m2+BkxDSriu4et3bExMwkRnWcyqAAXR9azBTgQNnestzw+VlH3RoREBmRpegEai3bq+7vX8Zg1G
C/ckcCIbTqbLmuD889SMaAxp+4P0hDaAtpcpl34htuqLDUflj6N8mofX9K0UO0D6Cb3JBiIaNga2
LI8kTq7RKDu5V+qCmsyDvyhOvNTSDDAMbQ1qKCm2MIw1z62trRBfTNn1zZfge/CCbLVaPLgDp/rv
OzcYW4UvA4mEC4S8nLNE5G4fYBy0x8lpUQV617TkhQ/fGfTilbn39GpNgh6jX+kfXXMs5al6lSyD
x/Ei7z4rJ52pDrxEFZiQNH1G4XoAXFxjsSD3UuwsqrttxG1QVmyTtCKaH349LlwE8Y6eOONOdKBA
8W66HTcB5pCqO7rU+iTuiEctEKcIR1JigGLn/GlKIvdO210l9pPtRuiztF5/A1E4WqtPZeE8l4DZ
gD1qJn1rO6PjTtsS8CPJrMZXJlXEfB6Bq3Y0BYc5UOSTMFP2Ng0YE3/HkQod6UIP1ksXUUh07u1+
E4yS6/SMcOzzZQKEy2y0O9vKKZvMHMuIejz6CSrPEWLlmaa1S8xBBesWPprY/INKHiixes6OAbMi
4RacGKQ6u7b6/EqKfUJ2+FyxS07yPuqthxmbYWf2hAFa6CKRAQQlK7efUnyxzotre0IAEcdX4Civ
CB2yCKmt5lK61kugYw2M1LeRuIq31HEFLnGbiSJjn5/Za54E/4DoUB4WUa9p7x4XGDShEe7SZa/y
KN9HUpGXu3RjBqfg42sPE5V7t2+9zci6us4IARTqjgZ6164Rhzn1PrfmvzE9yNCFH3lvu4rmS8V/
0oO6q3eknKk5v5YcSkejL6w/gVRKMtXie48q7rGqkaj+4Bu2TzoGLJqoKntBw341dLomdxHVsU7R
IQubYSqD3tsEjuuujoWBJVfmik8KNZV/FfZi80ZGc8zawMOXrrIukf8CggnKtXtXLBO/ac9DtLZm
Nb8O7OugPyIT5hI3bW/4bzv0SgYughhP3IBHAkSb72fYMODjQhS1DOI2flg3AkC8lPGdzleP1j4F
Lri5h0aJVX71Fkl6Ukk3CH3XD/ZgTaaJvC/sXIBc1VZNsNkMO+AT9XaEymBTc12Gl1Gr/Vhd6NWK
tWmBFAjjxaUJrsuiQt3jx8Y8+1zhPg3CBDaqhEgi1kPmWNTwlTRA7EoxFAlKd1nAZuJ/S7oegtnH
kBMjxEMvFDmZRfQlN9gorXYRYj/FwcoEULkjI7WLgIGtC/UVY85zTNpmbbOnHHImBR8VYpMYEJck
Np843iwf9s79NnM13dh6jeHPpTNnKUhBPrtgG4JHfBaz4SGNy2gY2q1Xoo7xhDiqv4yzEajR/Rzn
hOgjK9eWxaU8D7rrUf3NIKJ48Ng4Ji9ZEAZdaH5GtxmCuVNMNNL4LSLVHvr23VuLpRT1Px7Y1Zxy
orhAKWsF0kZyIr9FP/dR9MIb1T9KHiR1VChNg6xYrb8uaqK1hMqbwSP23cC9AiYzb5uXnisgPD88
pvEuCgTmDgxOsyXk3DvMjn3s4T4OeRmPOOfwfvMidR9yecqBZDDPGlrgPZpuNKbq0J0Gxbn29iEQ
cR7jLwpnvxLjYe4cSrgJh3iXcXF4rx2kV3Imtm3qD+XmLRsOrjdAnsG5JJ/C545gqceJPfzZUNsf
T4gNB82q050Nm4ZoJ9xb69yuWyJzkAD5e8fj1bOnpmZKTeyhP2oQhuxh76qRvVfzpVqJzCTnAmHs
5CKTHfgmpTea/cXmnonYkM9uUUxy0zA0brmkWOzk4D6CNHOX7PX26ZFBljz9VfA6iWYzHwMyxVt5
DvTSIxzsZVcURuZY/c/eGurfenC8kaDgJGKpe9mZ+PxVAkuGVP1RmU22UUDDU9TpFVZNBOj0XA7W
vmtE0oG2zvD8yT53BgdzxbWsbsPVgeyRG7Bi0djyVYAguW0vK9tvuM1YFUd5an8CqKTuAtKwexE/
YmwAXFoTtFNlJiCZOJoQn6hlam0sKQXZs3nASsGgW9W1JrAIPykLLwKS8foYPpq+qHlfVZJ2CCNm
3Wc2JIMPaHX5xPwpGbAvhK5jgggeiuA99hERO5SUWMGYQ/nS6QoQOoov0D6RWLUvnmHViJPeDqHK
16l+rev8X0sWZUlFKqdw332cXWoVsowi/Haae748w+V6Q5iSTU9tR62mFA3Vc4NiqudKUhekvm/B
/x7/XOLGiDt7mXnkcZBfrwcwU04L5xk0ioqQtfzAmv4V9/wkaSdmRkdUM5u8Im0bWxkNQ2C5tFhD
89OFKFsKMSi97CNM3BgGDmYccr85Kyha9R51+u+fhA/tRO5eSGJ9HKsv5212nBme5/dhT5u7UtQD
5FdxCfpkAlJksos6/zPxHQylzKiunjHnBgEX9yWznVJpRDBNJ9gCkUoWccZciTLb2w5l1aDAT8yC
IHa0xyruTAjqccnLufSE9qm2PGosycr83Z7UrqEHgV+XFRFY3SOgof20q1wmoccsQmyO4K1XK+yK
7tlb8g5EDU6q5EXI6G5o2ChscwzpPnQa/l17KabIrU1hxeaUPRF+cHG6cW5OtBgHByAosLCCDwjq
HrcYtqhR5uAAM1y2xy5Ui3jIsvq0cLjflh4AWZvnnYJWsAC+/0m/Z5Um3mPcZy4cEvHq1qpDwObb
+A18sSkdu0gS3LLHCEvMIkbzM/7caqZXCPLrLf8Zi65WWN5VMMIrIHo9YuhZxgTDtiKWgZ13rlSB
TE8XLuEGev9IaC0UvR3IKw1DiUdzcxlWB33ete2LrlyFV7ulNyADHjrMBTta0aEAaRX7uB1id2Ys
kRNyPaPEuBzIjy9snS3zvH9kNAlHtu4YQZhJegNavvE9VwuUuTvWidGgnFZL/TqzzU6foys8wDL3
Ujr52a3mYKHvuM6sBhJgGKspGxFFboAP/GALn4nVivMKtSLEG7+9BdrmnlBHxAKmiNdqnK+djlwl
WbrdkU12l9Jvu1dUORlbFStpRkG9y3RIWWjNktrdW80hpPB+Xlrz6t0h5t+yhcrOpu+NTsng/mP6
1HlB6XW7NkxMI9uBTNdnckF6LZDHn/ZwtU6YUF4WMPaipywxNQNQNyT1iBnkoicWHW1Xym7RiQ1R
AGWgJysnO4xJtkWS1bLZ8FdR1RMV8zuUUUnvqVRsIr0bKnqJuMgjHaLUKaGR/tr87pDkdGmUMGHA
RdBbmDCUv9VGyMskElpQjuACKt8QbMezLYIbOyXVHQp7t9d9JF0bBbmKHw4LZ2WZfmgzJCl2ZiNV
LbabJWe7NGCp7kZElbo1Q7/DIZkS1GY3KDJ/UjM2H9vJ7pylRGAKDT6ZSwc7lASHAXAOdjUCXhoE
kLJqdZHYaOSJ1EzrxaDV2gN3rm1dBtBuLDGKVewXk/e2AMnaAup6UEp1H0nVZQxfn7FRk1UBGPlQ
rbdwe76/SSqUn100YONgsvoySppWS6KTPsDj5XDo0JR8XKT9vRR4fvE33i3UZvnQrr2dL/vHijBQ
vcUYp9CcHw/QRucMptmVt1/XCe0QeqKdf1fX5qXdiXlUwzUP0uVTDCdsNwmAIOf4C6h+7bvcfGRL
REUpnTx/1poe+Xcn49QI7Cz0BGXLIfeNl/9NGj5xVqGs5Pw7kvaxEIgzZHCA3mk8j/wtxq777Y99
Y/omdFeyoS8tWle9ldR8RNxktJo5xkdu554KvDkKR70Wg88BaFWJ7cXgtmTjKGRGBcdnlQrXbaDq
rJQIgeuLSlXVCytVmqdA/sW4Bqj4UBXWD/kzmuCXFV5fX1Y69+b9Yl273jIbTlEaQYD6zniOmtDu
S8KGyKE4MzPS0ja14D4IQwJEGKGW1E6/Cd1uBx3D8Qn9mlTJx/JHozI55jLKnQ3lf1LYRWxOfSUX
HXrR6i4phqy8+nWchJCB0vQvy8X2otizwGWQsU2LLOuJabZKhOfYlit6RM2/fXr6UD1Xvp+aJOSC
mCGA0ZY75cJvLzv6BVDw1L9jXjzH3RRTFrREWQkckY5uYr5EFj82Uo2fDk9vpftXz93VQF4+pZvr
D2cDJFWTu7+ihn3j/4DFEpWnkYgwp34bCFMsIcppPM/c8k9DPqp1XHfKN2C9jGUdU11bGyl9Jmms
yaI/uXA5gAw3slChW5wlIfF/LEzMEEHNqtVGlO7SHUMZMHvl96bjJosiPh9wctEUaFvH1OeNZQWM
KsGuaYsJ1Gfdn0cjfTyhpn9yIh4BX+NmesK3D+D/Qhhc29a7cSdXJ/nZdwD9KnPbmzq14u5/L+uX
6NF4owKXJceqv9109oJXGO6idOytRiwiCRpcc8Qtd/PSFODyrBIpRsm+zNjaPqwc9oswEGIwUccJ
niETeeVzE1kNlZx/6dTfVe1aXeDr9WeGoXMjG9hcjrJlDudFYrVRui0nL3x/2nqGFd4oCEsTzCyS
wYHpaWgmA1nAx6uOi22XDo80C2S7HGqvrQixdKLMSP1pIVYkJt5jtIoA/t4Dio/tNuWHoU31vId/
Im511KPBmrxOaLzPwhF3w7xWEnTv8biGMHdPr/K5oFlAUhMc7I9J6STTpqJS/c6vHQwVMqxSaT/M
12l/YgUq6yNMMCzOROK2Bk6h47fEFuIfaFDJ9hxhb1TAiLE5y9aC2w0CjzyhR4ST7mxiTgIPhZwT
GKFZmedCDacf9tGIC0KvcenCwbVsbYfW2zxCxNBW3cP4B3VrsV0eFFkGme6reVScwpxIJbypNx8u
nm+ziTSvAosHq8jqWZ8oqagQcxjUGIabqeAcg8nEKH7I1v6QMk80lAnLUTjhyC1btTycgEBcbyEA
z9FPS6n8068eh+ZNDeDC9+RAJNCJX8Ss5Pm1YkApBEMt62EChaRYy2m8Z+hiPL94GyWXBskI9lP+
k8VS/d5adHeaAdEkF9HYhZUWHdO9zvvhbQ/MT1+uQ8QFKgn3bWqsaejmEEsBSOss6dkTQHDvtKv3
ASUf2HBrhi/XNIJDN7nvu8zbj/LWRdex4/l2/4udQ5mhd0EDEsBz0zSmtEMKUCLi1kFNTfcbJqRG
+PLOI06ZP4TY5sQhdWqKUBhZJbpRn97YBsDQ7km7ke5n+kzcKl8zXMLbFhJyUQqPFBrKS+0sQNxU
dJLnYFk+T8ggUNYKu9RUJGeO/hyV5e+OJh69QoITGl39SUzbClMLa/zEB8gFD9Efm7q60JxDvM3v
LaR+OZXYOhSjOblptoA8Ar/D+Qfx+5wUwTip+bZORQryMpZx9MVNml+CuZtMBwv1I7/PBXOZo1li
ZmReMl08YBaQcqr1areDLvF65EjfyKHWpCmmRvwfskBtPQl+VgrblGQR3OExrbvoiOQr9jJu2DXk
l5Jcc8bzwgKow7Xq5Z01UTHGLa2oHhJBUNOlW6UYMkfkk6NKwJN+74kZVgwBFD/7QBv5nOnWdP0Y
PFBeZTWhxefDCDLMJY1Xvt3iuO4ZVBID8bgFiMBwnFtTVsr5e48TpEY8o1K2VHu0caI4VPIeZ8L1
nqMT+y5fUq/o0i1HM3PnbcNXSvq963VRjYHvYWdDZgpm0QjDWt4huX+yaRY20DsY/49fQY8D5nXs
XQ9dq7daJtFXqWChAhn80DUq5e9xCOZ3j524WnMfrU0b79Xmtj7lj4AaPj4OXntilBvLLbHnkrm6
EsEg4gwP+VEFHTLomF8/E0OZy+lW4dO7fm8hVwpZGvVSG30Ma8pNIMV7JMs2xHmSd945CF1wDx/N
lK7STTe3EsUKEVv6WFqG6nYOlXVoCInsWMkLra2E1iDUA8EopRfpBS3zr71PpDiLULpr7jFZlAEo
I7d7/3oq5KL8ai1hU/qNpRiX1ednPHKHuDniTDrjKvRXaF6T4/z0NlImffFWZRy/B9QhLp2qr1s7
IyWCwshqE0S1g/nL2PL0DkqvDXOb+aVliLpKlw3+Zfvqwajsc/xDwFxW0ldkLyX2aAfqNOJHOVlR
ou1Yp0PH76ffnPGohoHjfPoEbYbTAyviqRd3bmD+VdEqbuXmP3XnzoPIkPbepYlJ0M7Va+dLUavf
UrD7X/+B5RfAFBE8hENhH6kU+mSx/aaJq9JMEF+DIy15fiBNADR5Ak3IHmdPik38cyn5y1NUkPyc
CRsv4bwcdFWRfhh/y3sOxaQs3dA9Z8iQdn5ajBYsjRq3pAxR7XSWtW+g+p5wC3+xxYsuVRNhYqZl
EeVo3aaE/tC6HN+XHoUZFEMm0YLY+BgkzpF+0dn08x+oTYbq5WIoXYl6WPdERF94/8OHCRk2OUGO
8Y88BH6td5hz8zDHR6xG7euS0LXZViI1x6K3hIWr065RaMplqkhb0XDR0l0st3QBpn9Y4pwbVTiJ
Ua4YH9CnEOobylluXeju5Vl3AfUAENRTthi5h/zvmA/L+QLt2/5VobJz0TthzCwgGLt+2AaNpYj7
LICk2ndCUlK4RuBBaOZmFp0OM09AOaGFjJ8uH9f6yONN5kAA2WiEGse4B7CVt5q0yEW1U9CbXbLM
f+XOviy2YnCj+eGvyNgBU3TyPg3WRnpd0eDXGeGyXMjCFxar/lAJ6Tp8bwGdNWiLN4hi129GUT4l
uGC1nDHq2AY7BRrq+J+Uf3m8ljLUTbf3JhgX3SBraC96uA7ixdt7/YxaXnSMUTdsp170MJMIaTxg
BYM/ylncgft5lxftkPAhlBRKKik3Xd/YcBAb+Q+e9PsDSUIrtAtBRSIelCCLhQRles5iJ1aIrwFw
ahphgrRaQshmN2vienprdNhokQNPu6XUoVEDRAsRIUpNzYqLEImCpZ3lYY2WqiKesYZBUOm/9b85
NQJ9XBqVY+8nwNrowMft2h3PTi9KOIEhn/o3QJLG7FEH7gSIj4/x1AA2Zi5DUoQYMg9sB0XJIqgo
LEg9jgIPyCnyT0H4PBoxAvG6iJgRjtZWUDwDJ4j1x340FUfiKkRtcufhcphiDob+5gp50No29Ou9
b/ES9DwjEz+X0BuSO4N4eDWpZg5FR6ocBSKZ0MqCFKSVnaLuzbdJd2sZ9mXjURFxZMFnho5uHGcA
mv82coXUnYOtgmh70T0YZN4/KdTgtNgV/7Tf1UTpGO0oKO9tl7YDTv9B6J+uDojxaQi8Qop+Waj3
pSX9B36Nj5gpvGCA3jFTg7BgbNvKeXo8eWUSCdWuWmN/HStsNnZB0GldBYCoomve0oLyNXXTQQT3
R5SlhXyVAWre5IQqblTRxqwqcgt53ek9vwmPDQ9UmuxE0y8cJiN4I0dKLAVLKlt2amgRgvy383x+
hpv6DdT8A45YLhNkQuhvWV4ZWeUccroX7zIVd1oAZ8X0X2qO8Inv0CELegrpyhT4LrRz0BelmCce
UXLmRGrQmabv2zgbrfmDaDXMHV5e/RRLqYwFuXtpqIjVwblhbIU+xkUeBjW6xDeSlkt6dYU2qmYX
RfGL33aoD/z/RB1UAgiFPeIA7s3UZL6/RlEShdhLFjzXOrmlphBAwkec4XtlhvXPAGpwEd9akagF
5UIqSG6gEKd6WbGYixYQjE1lyKkjA7Z51MyUWSRao+QKTKBSrRjaSMEuGghWEbxOeUy/vqU0s0s0
fJnUvUtJdGLanJe1uvZAPiE+Hh73zIA6MH7ZCjVlGP4zSuBYnyBA9HUX0co2I7BBHrEKrn6aT8cx
r9iSf4MFiUDyDzANhzw91wIFLkFa6Bvif7wwnZC0B8HycsUDB1kGaB3NXF9zaHPFSZ1QonoTdZB9
lhWFIPACrHm9tB32SE2R1i6/hAzcGcGTw9yiekKDaGY4B+AFnA5G7ZVeDsUWBqoqEC+Xxv1Ur7kz
zX3D+pPjQDAoqHy5S0QwSR+BHpHAt/070Z+p8/ymTan7EeC33N166hyL0YI00qrDDwKHd1h9yJZW
Yk5bxehNhGe4N9eNAQy684bwOeeb7gO4J/VUBiLN4Sa/gPslWZlmvIXSjX4pBh+8L5mdB4smvz5v
dXfZEPoU38yivk41arkMLsz6O9LPTe9gV9g5ykyH2v8bdvb2xjl0oE2ZXSC//rpdECcVKNYqnDtb
nMywyBNAnwqdid3nL2ETBSZBLUJ/UsAbZPzeuI3Af9pUHkqIgYB2bMUAxInmwb8AyLE6pZTs8E/5
dJy+2fsC4lxBcYs+KpH9Q4/XcKO2H4ShnW10QH8kZEk5XSK2XviTx+vGp5y851ywnrEdtTEUKRKH
yjYCh+wHWhKmSEe0GYwQBRH7x1cEFnSS5te0g/IrNmiHKq74pTlGP8iVxTZYCSM5kokNhBYKcdb5
IwLmFdh9vL32ChEdC8jN4uCb4SJJrrT6Vqn3w0YnJRwoX35lGroJ4HzUXguaGcwdsxk+NbHwM4y1
g8Cp9kKLYSDX1gf2UyTLxpD/BzSJc+byLl53JyTlH6YFzmu8nN1+JywCTvl3EK5UxAHKAyM3dqeo
GD6gJbq8qRxkajw3spkQOhZoEcuSi/4QdheGlbrCamq0tLsMBw0okLT6JTdv1Kky/qfaNLWkg5qH
9JcVnzv4rhr/cpu4xuazZXRWP0ixAXxKXyFp+lnZUbZlk1TSgPE6YuXuc6yws9HghHloajDsH4aC
ylnYDt4TlqZ1F1eZI5l/jvgO8xf8sHhHvSzFPL5ieADL/FauBNrtS19RuSymrX7rbOVnLaIVp7/D
/lyQim9k+jbQQjMBOgPLY0TnXiYYyUp0c0sBEKZE2AUNcsvr0iDfgn93K02H/H22OEdThJ/aaZkz
gvTNLYrOed3wyxv7Pp/XH6hjVfZk9xDXTyeL94eE6680jx/JJBHIcV8V/51a+PQ9O7B9QWb8hSd1
S+pmk2LNLkyv599+msGyKRJ9Ks58x9g04tJxPM5zyHFQBHcFo9WKt21lI4zNntUWOahFBc3PFX0A
+pT2jO1ER5NL6VA1TVKLBla3/Nv8gptzf8vCSRNUVqjFN+jeC1msiLQnPO8Rv0dD/KrMH0Qvtkvc
8/Sz4NxO3vmiU4wUTSmCeEWlGqs0++CuzXPQZhRi0L91RQe/k4NgX7uJsph3Ka8PGpbF0PpoJ6bX
gHMo1QIcLrIFBrBYg42T6jrJfAMJovbGg7rq/LcPBFOqMepeeAcr4ei9zTLsBplNHZeVFpqobtNJ
sAk8VKKbX6fk1lKsY8YLSHVvdy5Wteau9FlMr91ZR0yzuzqEp9I7QlvD6znVlPAS8Yzi35hHZF8F
9Yb4gcewKS3VpFTCK7h2CGUGMEOqQ136xSSPpR7POmBT9C0eEmxwHevOVE0ajHp74vRG0J1kCU5J
tVlbJkwBX2x34RS+xnXdarB0E734PO02TGItCH8PqXUAjnS3n0H7SEn7SqKM41TJu/Uqnk6m37Ec
okAqDcagMQOwbWqGbIZRVEnGjJKC0llkDA+4TSYMwHHhLCvzzx8BFJiV6A9GY5Z2ZP1WGeRORFyg
8Op1CEvslnRVjkOo9iJdAltzOlw1+th6wn57+Jk2pxp3FZuigeoSwENg6B3Ms7KolfrvK890N/3j
NfWKyoZ09eAlU5bs32ZO9D66WgWKb49E+3dxYT6AbN2DA6TMujMOTuNNUGruhrp8rvP6RaD+sPSY
tCJefQ/uTYmDhPMKnEvu5/FCI+VtKe3oM1oT+ttuAMeUnMS4R/Kt9quxJsA5siXXdTUP54X9RwJ+
VOw8oX4Vznuluf3z9AZdRt+oZw0NlPxx2b8x2b40u5WJnAGkpqNt+DKHjRNSRD2+I1Y/20oCEXIJ
X/9qgtEh4z4J3h7jK7kcVCNY9eOEMz/Xj4mmk8U05gGh2bsmJtMWPBXD+YIMpeKXceQgQc4HfTx7
sqzU60ryoG09P3rFMs/2jLs8NFysFsTbWfuPrkvOLEujZu3CJrnUEVWCyc+SX6z4mFhEMT3kFj1o
NQBoqrfHlm3Eq2bL4X7tirG33GFtRKJCKs1Ay1Ikpxw+/DPdx5LFJCRxX2KCz1ncwc9iU2XRakck
9AAY2uR8JBWK0StsJhXriPh1pA/4P3X5qjzVcxuIV1Uaa6KCKQJ6GxxgUUbhmfg6qAPoNreb74un
0Q4a8GwdyszTlyTmsofL+9aCJs/J2eEJcOHIM5bCT2UHkis05hxy6+M/dK+feQuFOnKsEWbVH6bQ
WB0BKBg1bHCpQBF6mrR2O1fgZlRtYkQh0vHqevJ+wHbRdk3+FwTEhfIqwTPvrew5fAasE6pkkRHV
ymbaP2egWQDRKR/0ge6mXNvux1qMw/nBVhH1vV7XWub2qyHq/3MYcTrO+AOmTgQ7w3enhppdkzAf
SerrSTcNbjteXfVhxL2A+8s2VNxcN+5HexkudZYXVKM1hfPRXlnLIcbmukmgAzIcS9wRjEurYHMR
Ar4jNUpWdwEOBEf/6hXSbTBTPCzO4y16I+DCPANH2xz0lThaSO1QCEz5TSIXFhr/Dz53Px+JT/Xu
GsLA2UBZRWh5amULcY+nsZ3btPO+wyTbPgKtX/eAUvNWzs7Eomc6a/uC4Ozwdc552ynBcg6hZ6QN
xPqa1psdIBVX/q7CV2Uc/TACKixwMYRT1IqrGcqoVUVj6pFYSxMnKZKdAMYfON4QEvL4rcALUXZP
d42hB+1Ga078REYzKE5O4qO8/wWTki2qpEoBEnAqT3YfbP5ZNwB3FaBEBGxcpGN0f/EOy//lLmIE
v/0OL1rwkKuI92ta5g1Q6VtI01RAzafdufmRW2sUUPTT2gLC6g2cgcWt73c/712fnRTMPLFcm8ae
f5BEApTq57jlJmbEjnqH9hqitDwxFklYQPjHT6Xy6cG5kkEXhguOVortx3DJzw75HTGFuQ707KBR
lMzbFQt4HuL7Ec3NcKtD1KKDD4n4tToMP6lZ0cdiBhxDoR+5vit6hrUOEwT0+ENKeaU2cqHr17m2
hzrSmxyVzLx87sIejeLXp9sQm5P05Ml53gf9GGVY+SWfJVc4bIXNOUwbGpUW8GgIUew3M8yQ7Suu
pX07ZRY5uRddj7ZWvO8LLH5wi85XRc/uoiuVDYB/X3FeJyn5+rs/rGuPbGLjD0mwKiHRS+fqXf+s
35mzDsXwc7pLOI4oPJ1IgApVjcRxevJx3YRHMkqNsRUal9BrGWIoHUx8gFGHJlxJBAmDwm4uF/pI
dHbaVVaM0EfV5YvrSFLp6vtS5A7L+NppLBEJrUUGs2PuAdRZR3+iCLZqoTmDcVE+lOMGAGnAn9ss
sz+Sx2xI80c3ar5FsYaMmaYqy8xAKheLb5E9U4YqKQMR11c9qI7R3vtAtFq9wJaqqFCozceqMjmb
nsrmljxb8yrF3NqSiQkAs7G+o6rL4SRvUegFEZYPUX5nnh0NfTbMKlfkZh89XKcFFq/1/v7ETaTZ
kwJ9ZOatzw7VigbBYgRHhWcgClgNRNq2uD+qvQf/4ZpJ9qQOZdTx1F5SOqSZAnuz7tGFTqbxduTt
+qc7fmsKGuZ/OpE8z8G237rvzUJ7MsLreWn6sCvrQCrepR2sQrq5CTmsf8A3Ifo+d7oJY8tjCYlH
8srQZPcQMphnqaDr8jF9PQVca/nMOsq40FMRZLjTcvBFfH6GxK3ZJhp1+WUH5VO1n/Sm1Pwo9aI+
k9kH6o0PbhExMWF0ik3YVaG++moOrlFXRFiUfP8XNPWHovVn3aIOWtYUbRvVAmbAClxv4tLxEb+o
mNkOgput8JST5u7iazLnVa+dmXmdaR+TXM/WJ7DCHORrTPJyuZz7aw2XtmDf/Cqqx39O1zMFMGI1
wxamo+9FgtgmueZqSJLqD3QpuFUiQuW8AHLksseki1fOCIyDIB1c77xLRr3EXuoZcW8+HuTWwDqW
sq2Nvzp0332Ozsn35hZpsV69uTZbOzPOlarRTGk/Xr8Ni4GSpMHcSFAyY0CvCMon2Ysg6uYgkaSe
jVLYTvg0N+ZrNX66zxsehoI3HyIClHC+GZ4Z5Xcd41kfwDc8x3AixLePNANFXcp4twcJ+lTtjkoV
QnmO/SGxGi2xyBBN5TxmuXamsjcFaQe1hBloaIxSe72YgLLICcNnB24JipHQ3tJ8QgUT60JoZpL1
LqYBWLV7aP7Y45fJ9xArWlqnqeuWrGKCgxuM/jwZKWeyEs7V5cUrU2cc/i0m97SmbRi08HER/600
86LOlyIboRhSZvNvo7bZHh6n0ZMxGAAx84nM+OBcw3VxEsSc1IhkDqQFMnlIUm//CZONNABxRIv2
a2YyfU7QfmO+eAyxzjv/1hUUTpZ9dF2n2cjI23wqtjEHBJWvIShzEjLbhWGifVlE9PUnCGiBQO2u
LiglqRtXejzOksnkh2jjXPRPA0vClYVjeSKUPdF7XJHmEZ1E4RHgt7NPsbra+4+28w9Wj5/z/JiY
1K3hdJRaAknRtHdDcSexzgIsWeAqrmEf8w0LNgr8Llx1a+PaAkfSfZmCUydKtmDCgXcXxCAw0iw8
t1cjLSz1FFedwPDCwiYChi8dlOJL7s3t6YbUl1fSVzfomC6586EohWkHGx/aZ3xmVdR1reT5QKmV
oRlNFFWz8E+KiPbyNOGa9Nxe1NYZmCFDj4VUIPcsoBr9HSBUNvmIagGN5l2mYQ2z37U+6t6P9KnD
q/xFJVvZvi+AsIn23X24re1LWK9qeQBEcmRVuRXW7aWfB16xI7iA0RLDlyp+tNQ5mX9qiVohPa69
A24s/mHG2gICYw0JTjh7Txm3WfEnrN+vqS/L9pca8OWmaqcwVPRkdwN0lJ1/sXfXjx/oeVPdz4DT
zjczCqsNiaqotqsL2JPrg81t5bUa8rdNCQDqBXQamkrDtCHI5kmtqvNHIU+dLUBrMgZusEuJftlZ
H0koP+Zx3NDm+4z6yG65T9/FwZK7J7Jm9LxBU3q7diKVZ7PYHu4TvPN00yNuPK4PYJTvFXyqe72r
eLqVANwl0KYHU+G6fzKlUn5H1czypQcucWbY/phoVzp3e2mBwW5PXe8/ifwYdnHlnGXvovA2nrhw
FIlZmCLYc2D4NPY0iDO1URpBjXNWSA255nH3Q7VHTyEMdvCZiWC/tSChPWl9Ux64gjmD75psxwBs
41Ln7149WvLvV2KeOH1buVnqYbfIBlYM+J7V2ioK+JOFCyZVqnNeTX3aBnq6CzLFw3dFizCpS3rj
lF86zQNUwBRN40uLd0LW5sCuVaBlDWlVXRxYcU2hXjdgiydxHf0K0By8AIbEmIbH1Z1i8LkSdk5V
a1MYrzAhYzEGRtaCF2F7keGnd2Ya8ybRU+ldy6IFJHnaJBx1GuBZTYX+uBjZ6yX7Gb/hDZsiCVj+
KAD5e5kHxMuKAF4jO73R45qz1ogwPF4R3iSVU16On/PXqFS3O6DRAHzHni9XWbKyxoWEeeY73234
p7AwNM8WqVipVIHdNSaeEXIdZL2qrezx4T7Q7PrSxsiiv7p2GowJCm52xSIIEjZH8O39p+ZT165G
R0hm+nshACtcs+YEEiMiUYHXqYvYl4ZcMq87b02Or+Fr1CHHNgOYTIOZMsO30AjzEOb+D+qY1sUg
X8Wk4GC9Z9DUDRRVo6HC6RiP4tM38i8Vb9w6gT2DqFE+3c2iy0FIBHUSXbQEldrk0DrKS2MCXvK+
1XNi5HLTtjEF04LjyED0UJeS+3fV2jogNHk8u4IzzFILSp/xygH0ZHI4xJ10DVS02as/MlOeY8HI
bgx9db2kxcySm7X7KkmTBx95Z4SOvsdqDNJjeVTRk4HDLX0u/68FDymi7dOQURHA9W5gYcuSQvNM
9oShfoZe/siE1tfneM7X/z5VuiCDuybXlEm36b2Vd/LTQhiPmR0KvlWJ1PSOujiNWMphHxBg5cUe
xBeiJlWbKj3qmma66u7bjOEEYUwFP0FwAsBjMxlItBV4mc8Hx/x5UmcNOXkraI1ZVDv9/17fL6ef
PDHZzj3GfDpme+8RCnRV1WZz+H3UdR6TKfvnKH0CblmGua5rWnxaTtM7QG+iEbqV3z7rX+KGiDuD
izx0WWWs+czy82VqqkXHXxkXZYXEETL1OVvVb5PAJgf56XmiWjg1JPNVhxUJlSAXh2pZTY2FNIZd
603cgEENtINRkhZHiz934KudFtDVA99YrEQgeHnYeTMKXMEX9HesqISFdUFCLUz6s+bScKyiSqnx
G0T6YI44A661Bqxhz/a7WCrC0SCYo15gOG0jdU/f4NSWGz4BRlnMAtE+YC4AWpO3u7fRvBQuW3h9
QWeNZUysk3nrxcKuSGKNj8u+J2MOTOEq8Ebq35AGjgDLINzhiauHgppUgTzz/Cf6ueuGGNWONjV0
d6HT74AC/I8KemBqfrKPpxzx3KxL/NrycNmXxQswtZNG0BWCJwnqkkIHTg7GMxSnNyCnYwNvRGpP
t6rDKyvRSaZ28uw9S3y8uBap/y/2vm+9CiJxmULRV+c1cPErnE9V2bkPlapfOUopkTaT7NAFG0jO
qpcOFaGDKh9uxDDOZyCMn6pckBAEBNIEw1NZaDkmzfRYwrCKaaFxUBxq9PV+ENy6THbPGJ4zh9/S
+fTgDrLdE2cYz5fWLoQizl7av7dMe6dc1/D7zRxLDd05yIshFdJdckYs+RmOGGK4IzSib1s+XS4S
1UCfAAbSLBeqOAQFBAPf18o+/M6h2mymVoTjsG+VMLRVrpKkmhjCLzPg4rd2UTi79AdrxbrKIHgY
qKqVJd93PqQ9XBpMgle00FwWaLgkn9yq8MyHXcVice/M7TLURUfwlgQLStqNCt3n4zRQ1tSckKiy
BuudnweGecnmQMMtA2RgYLjG/zcaGlEN4+zmtZ3qIEpTX8NZHWPXA5S5IA9SDwNkwqcWUuJ7Gr5e
ZR6aldrBMlFgZ5BKqVrpUTuzKPr0s2sLC8toVuTG1AdFvT3PDQoD4kkC8GXVPBG87E6duROcZQtI
Ovzacyo7b9gBmd4LuQDbYsg9hHmDmpngJbmPFr5rgiycWEMiPZa66SyfTLWPBQ31ZBtayw9oE1pb
Gr/rip0CB+yPzJhRMMtPZPxMQWP78d3D6yrHMQ7Qjf66JR/dcT0/kuTmMk5OA76AkacyaQI1aSuZ
tJuL7wvWUmunhAvGFtL/NTzcUzB3MhyY8Zkhp8mrsrq6kOiZS4xcLZ9W+ftuLMfMK9uSA1ZOaN+g
hy1kOPo0MpTJviADOxVS3mSpr/3cS5ZFDwcSh+iDYM6p3zA8LqBPWL+GgRFP9IdiIIyR79jDa5Jm
8E4+D90GBec9P7eS2a4msP1nGZL2IJnJ7Edl9b7xLDLnkPhjPX17lkz0Yd3YQYXME6esdzv1Bx/R
1lyPDivLETFt7JV5LXjqUxMaTUKv8Msr4eEn1UXKfefb8UWvosx5oFDEC2bc3hYdeqQ3m2WA+L2H
KnLzGbCu6cyWJVwu4lEQGgpbwfFgmrJuDbndtXyK9BZWuuZOtk0Ttq6sUHePRZEbJYM6kpHsOFBc
LuELWS5dKzoqsUijBARcb94JagwNMKfjQ6/bGhzRBu5ajZLlkw4X4T1LxDrB2hntU19A28w5CEG8
G+taxYqA7kTR9nyywPNgizDkn2YMV8+kf9f5nF2lVrmdNw8SPNWjXSvQW88w5ikwBj3pCZKQvpx6
5sPWFO6PFcofgitQeq3n07FCdip3WImBoR8t1uHeX6Ww+Ly0O3XwDkvMOkiy+eGJljki4sMHlPrl
Ifbs767in5fPlXqr1HoikM5v2UaYi8uIxcL1ry1I2WrUSZQ76ksup56nfr91XHNUqOKPQNMSKFVq
bFMCekqNpbVCxw8rpYvqeCwk6koOeKRkGkXmmEJF3QMwidkd2GrnnRTjUlZdO9b4/PX0p+ZjNkiL
lQ1ZdF8MRNQkDOZDo13FegEi9pyFprdOaGziJyPDWUTPnRJAUQ8DrbDA2TZxhpfD5eGmeWcdG6ky
UC+GKxYPsbK3PL+7Gee9wbQ96n00QbuUxBy71dEnEuXGe6VK+yQeWblWybXXjBIJGI2hS54RjtYR
R9t9QvibdntmELQKMjiim0bI1iKVKOkiX1XDdbKs3txvui5oN/lAxEEqRLN+MBqtii/LlfXfq6NX
j136JgWEtH63CMoKnwoo7kRlSbi7kLuMWb1gAea30rKl3QCzDEAMhfqeYYE7KOvQrAzBuiUzAkrZ
5NIBDnA7PTbFXDJ08cu1mTKvtGA1m3V7wgP1zCGPpPe/mVynmHpGobIItpY+AipYEUJpm/pfSJS1
8FrQ85KL4vbG/ZXfhZoM5XaXFz0kvNF0bt4eXZjPuYXpnfvpSWEE859YcZkZ7GZ5ZQnenDIUAknx
2ZCzFc7zIi8UkQOc0vJQyjvjBoUk0iJ/AOiGMKUIAW2wZWCNAOor7VWLhkQoU9OwZmZ/+9FERami
w++/1a1utC6YVDOkKxMU4Z2kXnH24B3uWaW31eoRCg+74LtvTRRCdbyMHM8TL+nY1kFjShAIsMur
5d2i6hVbGlWnXZDWwtw0eQl3p/3uHa3Vbnwu595sPjEc+QryacsDTv6KGu79I//qFrjM/1f+SaUX
cjB3i8qHk/K61rpgoWxZlzUF+i1pAgrwnUKnbIyAyJ+Iue85KUHJq/ye0GyAPyjS5cZFWuwunLa+
wey/WaAXCByfXe+iFnizyLsxOayzOZmBF6YaR7TWujUaQ2WbfaULKpYz2schCuJFfVkufn0d5TFk
UflzFSbE3jvXwunn2M2Nk/Y6iAbII44wFCBpTUJzj+p7u9KuKWL1/wLtjWsrGNEBxzhccxlLDSjT
crEWi4jrv0uMmmAfpx5cqmrqdhQ/dkMU3E2vqDNxkeOmwBZNhYEYEYB4pycbwEor6eXICqvKs9x8
waJ1Nq9xdEIDhAiyqVoKSdMiSt54avhMhgK+Un785VHvLnT9wcHQtU4wcNO2jiO6ZRU1JXOpKSwG
SLQqr+ofUl1OL0Fvlpk8QM/Wo9pRWxG/V4Waqhn5BKQdtcdIRjd7HDzfKP33WP1klIy7yfLbVGC3
1xHrIaQdcPp31jddO6ZvQNhc8Al+XPFWdTfJVwZTrI8b1iBtoi93iBcfw+dFM6Ljwivzi0QaH/IV
CFMxB7gWJ+hI5FWmUegS5e9QWA/1fcHC/jJySj//pfDbcfsu+nwhi48UYnvHHLM07OGsVC781+kZ
O1GetHxrd+nsq1Ymwv8z0FgoDzBF8gCVtT/XTfp0YVOTuNB+s3xjI2cQtQ1f8t5NmjC6E3HXAIMn
mAxnY60xRusuiE+6fWFlQWB3lxsl7/UEUhMFx7sgDa9c7Mfdyr5zr79ow6BRvGt5UmSr2sUhVR7s
E1zymZOA5snWD+toyXWymz99CZhLBh73wujIXr0PhYNAnAjuEU5ETvPxa7VW6vnElSEqXeToDiEs
zuIUYwVOgX6ABPL34cH4rnPymRpUbI3w/UN3cKaoEddLeRX9u3ftmGOunh/eajq34h+9IrfPVBow
l1bzKkSRka4phBFTa8vT5NBffJUSZ3MEu6AgPZ5ZcMX8rDY74zVRidHxvlTaWELxj4Lox6UzX8Nv
PIIB6ofd2ab07xvmFMWzdicio88DoRnjYOwmBS6XGsoFsb3seX53amxzgyHdHPM6i/ZC9VQqb4/6
kzSPtM7wARh+4c81LZJNLQRyZ7Zn9Ej/RKS3P4r/j9fYKHZfTd64U1aZFB++yI/vmwiCtun0P57R
7l7A1Vxw2LXnNLJH1F4OUYXO0VoxctigEiI2LB3N92akF3P2FOGNQZrv3XrFJ5WJ62p4H/tNwzGs
0vDXNAenXfdy5+jvPJ2K+2t1MYp0nqBHTww5ftus3KyMHhEvHWwMYeevsBMs1/J3J0PiYeaqi6lp
3Z8KhtIgbvs9uxM16OagPGgxYBLbpY24vE2PLmOqAVCouqVyzovJix4JnYYVA4Pfs3P6rVJ3sb/6
mzo7yGIS/L379829WywVciIOSSB45FLVfPOhhFNHMpp5Y4lIAAd1vCRJiHv3FhO5SShpnbKn28A5
5zBcrIxPeUie6r6VNWHhI5cFm/HxEduWiL4o1XCfUS2dhUGHma4CusziNhr0CcvnFQSsQRnil3KY
f+N2lhswzuvFDuA5TDOSvI1MXw12/UzcjAWrp/5AOxduEgIYxCuLC4oAiOi78W5SRWY9spQE6Ujm
bDaID5HbCwPLD/q2bDq8wazSajfxDRq6uDaXxPqE7vB8+HQHkvlRqZfODVq5i6QKnIsk0S1Ad/Jj
QrBIQ+Mtg9fcqUFY7cBK1GIkpI1KDvuSL3EbCQ7/wh5KL378flF00IcNsI8UPqs9MPRquLaMN/w9
6k4CAoPxTS+6U2xousCvQEkWK6Tq4Lrv715cnrt0JczZWjbQEj3AmFuOxgwn9b3WRkiD1SwfOC5K
6qyG1AoMGN1XdlvkvsFfCBB1jcCdfbevJaX59b3TABka/5qMuwtECNkxlJXJ/kmXXJA4ybAFYsLE
VoMIxAVut0t4H5I0TLyuz1aujOyDiXAXydcqAHHjOy4kpAuyK0eP0RI7sc0jOREfwPppu5rOMWoE
Pd9i/unEr/2RJrZpKVxYlIBKISYRWINSNN8S0VBcqSmga1bQE+4n3EmhvHgu3Si7fsJFEDRP4US0
bOtfpKYtP9Ufmzyct3zBnUuUY97jMFF05qaWy1dDaLN4txkU3JBc2hDFqlahzGkutE0cMpJIYX1j
MAbPa0m5DmlnIeWGmgPA/+B1C4lbbmR26uoHkrXdzEiqikIMkvKO7yAvhrRpBIHkQ5z1F5Fw0Hn7
xC/O65Fnxv+srwDCTEqVYOfeMNtLOLF4CZTngbT4xG5eqJEofoFi/bZbW1zQD4C34mm28dVJZWiv
vLRjTLPddneRQ7mlB6aDt7dBeq+jBX6mZ6u+0t9v49Jg55ru21RcfBT8iEtVonp8TV4oOf+l3rfj
d7Khy7JuqDhHQMHKW6QCK24RSS5R4uAhdEQQbaSpgc0j6WA/7wpkrcQGKdf7PrL95cUQQTsL8kW3
xgT07EIESHM4W7FoaOOziNfQV61tMjmzSy6IivjNqiUN/pgpcRkuxQ9QOHd6gDhzmoP6ifwJGvD3
bwRaUQw9bJmYy/rVcJvQgaVlt+SMpgGRqA72nYEPXdD+p+/bpZsS4y2wd3o98wBB/jAecRCZV6we
iqRxZsE1/ln2S0KztWUBk8WGvDQc48MY/Tftl4/qmpnM3oPrS4ugDvXao6P2IG11m1NUlezepWgx
bMlOZ2F0y8oPGeV3/z1WZbm2inEuQXWapQoxmVc0ghq2i99dn9oZRJ5iYyj7IGM7I4fuxJC2M/FB
jAs2xw/2xTpmoDtOPxm9rOfijxP+fwh/Qza8p56ScaBSng5/PngiCIpteYscsR/xYa3qi9AcrBVt
cC3JOZLqOYZACj7DGgWQAIujGbNp3kWr4BaDyw9XauMHFa2sg7pb7b+rqFG1iLMvhY2GTVD7NBoD
xCPCHDGqKBCFG7H3D+tnrnBfw0Rsa4Qumy1yv7/9uN2Kr0PCub5vJ0fkFYOpoZ8laC2DCxz/+jPR
OUmAnS32Sx3ka4cs9twcv98u4ZQK6MDl2YDNQPzgt7a0ZYsox5N7oFmI2COs7C0dCbZrlB91w7H6
g4QcAFH6LIYNo6YDeicx5eA2oVGMZMVZrDw+xjcXIrBfF6xHmaVDPyewMMcJWViFXPp25Vf3aG6j
hZ45CCYMryV9m1BaUYWaads8A52t23TmymFJfQDXGikCgICOyEjpzHDKXhRALRcRfRhYAav0UbBf
67l0Z+qs3PlFERKftRNU4vZK+g6O+k4K7/hMznUFbqbVSB4B05577cC7GLNSVZvSP6l9DRyMSzLA
ay6xyRKTnvDMaImBL3EHe8A+YqPw0TMqK3BDbBT6bT27FQtXkwPUs6qF634oBUYNY5YwmlTrxu32
BuWIhDQ10ijgdOpnNafQwSN/C4qqKF7wCIqWvgTLlXpcn7UsKf8naQphL4JLznMGDudqDq21mRHW
jdmZLjWE0j9q+kUQcq/HiBcRvpJhIQ6xrs8oigLLqZl959jwEQTwVpWc5stkpDCMpOmUU1/vUgse
k7sbpT/TDZPWU2AaT9xAayWF4iE4Bd2Jg5HxxJlck1apLwKahVy5CcYEIm3xIxrNGnAixDSVoa6S
HMUUjrTIlyRIx06IIxE94aWjLI9n5BHrqhn6IIjI9ikhsMRyX33KTJIpPvj/3w7RfalZb+Qxymp1
Zfag5e86c+jCq63bv5K9er22ESU+YYrYI6tObJivSNbbqcVITXyPozqP/tGj6cUt9RCts+Hd3etj
oHUOiR0q7357KaCnL9j6c/IlW6DkBjdf1Dnrv9hmrbX8dcM5gtWg9G7vXt749QTCLX8RodzI9+QW
fwGE3j7TfKU7GsfYITHjDm5cMFV96KZDWnXrZ8TWPHTcqw8y7aFMBIwQ411QSrdiIbW3qpZUZuGp
k2VryTRhV3DqWI1k200CfZBEZVox7/0Fc97copRWszT/1iZIBi3CSzuN8bPAp22imRfsB85XR4U8
9MGqIhav9J2rYD/v/SXw6AFHjPmmwc1vFHDmdXeYY9NUd+fFt/xHV//ndmxqPJ9B75MBmgQXUXZf
8FgZCUV3YMSj/i3KgNC6bIK/OyTa4/zNKWxpBsFrRh6uCjBd7KWSqZ9cIUjGpy0H6cYgVRD7Ptfq
8FiXJSlfNTkMCwWoVCRsfkytbNGE0VsWF+sNCVtVvio7+Q60FhbxyumHhdRes2Fl1gAfv5A+pRdm
ouktPaDd6uLq6993gst8zspgiN4eKxlUxaktbd2ZpIyufx5Z620Q9GUbVLq7SAw3b1oVZ/OyzeJp
N3NNbEWSHN5iFJPykvTjMEvc6r4/4HEdK/ey4p+FeG9h/KxO2ZnucMSiuit8BPFVrVI1R4zwU36B
XkMEMNTwcKliHFCcIQBKlWaURXOZK2aUs7tdJCL+xcL3az8z3aVrcyVYTJHw5yYwY5Puqb9QLlWJ
QwZCWkqa0khts63zZnXYAYHtvCBJsP88Q2eqCARbV7m5q85XdQGVGPGrqqKCKQnxgs0q27GRqjaN
BT4aQKrFsilQoAOQAI2IhUfWATtUhffjXsgd9XSQy+YAmfe3oCzzcu0Tt82OnDceN47GjH7tN2Ow
5KwRCvzJYftsRkneSBoI9oXgyGSkdGsVo2t3qElDgK8JKGz4xINfWfsqYZV6jUJDVsSN8+99oCnf
PBJgnyFTxEmo09cZEVFRncUG7gqoXRDfFQQoMat6bsrFz36dPSp0TCuuoO+LarT6OzLe8fkBz5aq
T/aFf3XKOvf29uXVkEx8W32lghGxNVegRKb4p/1+yzHtqlX6Rg4t1cV43mwTF7aemVwdObrqQfWR
T1N7TMwt4Mh/vFZoXIr2z4tv9Vbc8Rpzfs1K0rp9LM6YM2buOs7FmQYJEwWzNRAb7phUsgyWg/2T
cM3M46x9N1AMW4rdtom/1/jYZOC+JCg8fJ97LfeiLwaVm6fqVj9985K2v3Gyp52FVSxV+2nZ/R+i
fIGNs2ac45bUlwv56SqXT7vY7lQqliSoLDsm92BpF4Hifu+rm5ua1O8m0vwfhznfLXGIUIDy9n1x
mkl1LA9s2BjvOP8FUqR9lvKu4cewpzXMPcjcBaMAnVmEqRBas2rdFsr+7KmqGnbhfNQ7yzx3z2Ij
HHl+L/9iqwxxkqdby+nO3VbU45dHJ6UpEtuMZNCjt2/0xqk2iQ9V73sq1lT2G/TUSIJJcwgaCwNb
IkYUDlJf017y9gkW6yFhUxbazmFMu2tkUQFudOJ84ZPGfMH6YDSyxlIFRjjgkl8UnHoH4IWh/VOn
uTj9RLgSXS4mSzyGPS7tayKv9w7pWRCckuqsNcoGltw5NcYJrth/yEJUlfdNTgpYSloL9KaPrM+D
3sW6UjdR05FMA9kDF97yLLUznfOLIB5wAu0YT4G1sxQqHiEH1mcTrZ9ADCzmSuHZbNplOd2gwYxl
uP48pe6Litt+n8Q7VmfZPhA6z7bZb92G7EMq7P4MdVFNKuShYRqBkzxbgG8JJVp5nmH9M353RQvG
NCkHwk4x3X35ZLzZrxYPO9BuQW6YujVJWjrgM7n1ssPfwlbuJ3YMLv9dWGcnLn3NAMaOs91F07V/
7ucrhcDU6u7zFgNm+MI9+RLjD7sJqeyflMZ/r9MvEda6P4KnklK9dxVSxSHNYeIPQRS/alBHVqmn
549mY8Cw+TSkKYvAs73KbkivDbjcKw/a7tNr4j46NxmRWB9Ue1smgTE2xh8JLkSxn89pgCoFQegE
MO49C+pgh+hMcpv2FGAh1U2fsn1ioYzBId9uYgA7O+io2gVEYH6KcdVzaecb+I5RTbzh0As9nUq2
UhKciT6BYFbnGmcYrp3TGbupFgQGnrJow3DTWy/pO/pBG6uCYq9c/QAbmQ2+YtcWG5hkye65Z+bR
YShwsMW8T+qDLE1UO8HeEtTG786Dkiw5rGPUxUX96W2rEYyFHlHOLGIwsThcxA2r2xAVkF//caQl
AEjj2CXMVyBBtB3cW32xkfZ0NYROigVgnDeeKaQ0MUzFH4LoA+sJogtZXOcGXniPI5AG9sa00i2y
8POmTxCnwhbKmugUxl1P6bcBxR8rvJMdyrEdNOaAaIJpI9SHs9O5OamE3VpaHAx2EAa6aGnJS7TW
MlNVgt6Ivq8prefJb7g6gu7nTFhU85r+fu16qE+F1IsjIwubZHLNI2x4fqA9MkrP+QS+W9WUjvRp
h3kxzBZ41ERk1xNmbYjaQAQZ2Iy7AJXtLvydr6h77DfVOu0Q0vDALNjYweMK4EA9EPKwU9VnTzum
vNyV0UVC9fK5FlzKxP6kJFXz8OOv8pM9bAnk+LyhkCALPgC79LAZ0JoK99dpqmpFTt8UIA92+ZN7
DoHNtg4RPrPrz0BkbRJ2m0Lq5Unq6ZEHdn69ckPInDh1qh1JMdavVc8n5EMlAOF6DQOzefCHjWCc
WqrFTtVvBlN/YnCc0oJf3cObqSXuv0RIVop31qf2G2iZGPtHLQx9WwMGsq6zc7xfd3FELTDkdQ10
1D4m70agNfbJ+abIoB7XK76Y+Z6Ko/fLPo/VXt0YRhmuVsh2Tgd1od6elnuSzsgTJC7wbIEytkhM
rr490iuOiyyObcgVK5LMUOHsgLZa2UEzDa5QivRXmzcbdldky1IlvC4L2H5h5rEN3GWYjPnKrw2D
ok8C9yaZY7wt4bSQJakLKF4oAAVCiabvZRAh1vvH8GcKnDNl0ri7PW+aIdn04LBBgnjww3uheLBw
0Y+DA/KDHqZ4Rac8x5d8QTr0yV9FQPGNDHyR09K3RQd2OzgP23bvAjm3HKqNSlUWM9heqvpwSWsB
nrD8P/qi0nTeZSavDz0xs148C9FL1LqKV2yU74br3pYqwB/R79C77lz9LeH2Uw5iY7UBjnenXw3n
Pp1Q7h2IjfCs5e5di0V3VFIy6mQn7qubqUIX+TKC2cYE7/CImpIhCXbNNkD3rkTZl5HJxxqtfWen
QeKaohvgv1DdedeAHeRZ7LyBD8Y0DdbpeWt+27b0S3I6ErOBZGIyDkUE5fZPEt2/c254qnWO/2At
ZgqVe4N8BdT2xNpOHYviqa6V0JgCEGt1RSkev9v9kEYDuw9SpF2urpk00LaNyZ4TE8Ek4chgMe6+
T7F1o7vt5UI6lOeWSvpwET7xFxwbWvqbaM2t8idWT2U50tJrUEMNFSqkZWZ1gIXaFQ4w7QjzJSZk
poXwLIoC6mBXszwPEeLGoUSYwM9Dg/d+QRLGAcrRBkfIGSBRRYa4snHp2uzgU6MgSm/SzoUze19/
Cl6jmnWDbNJslxzaZ+9UrhXk2SDeh39ykMDaIkEE7wt11lzPNf2QD3woBRLyy/3GPT4Lvmn/syyf
mklC9TXZjZNYOcn9pGb+dVRJQnOzGZiBoJKXrNYE72EnfnmuR66WIUc8ujrERjaZ5PA1h5vWEHny
9tRxSxwEEwimh4VZ/I13mRL7dt8EfFLGP/VQV4wk6t7Z29p43mMQv+COD5NnrHMw3v+iKyOk+DkZ
UoDQC2897QwedTpaEqQIdWfEI+CAkCCg5pSeoAX3Ql8YG9hsAEuWHt8fqSegmaG+aFFrKVityeaZ
nSubHgjUlFkhgmgE0bQ2PU1TBfTHseUUMN3QTxe/D12AG+TMrblq5wYF5CVttVetngpCBOhT0R8d
cWDGhMsKmXo/uQWGkQzBHHr2Q+BWy3or35I8tfGYzDUA5ngF1Z+9OEQAS2GIHa41akEEFONOSSut
8krEwAgrmp9VFsI8OGwQeLpYXrW2p+9PyrAEXy2jXblzCO52jQc8LrEJvTX0q2jy6Wz60zj1jEOi
Wm4eNtM4QtMTd/zqAbeLmxcwUc78Iw+HoBew2X2oC1YG4koQw4ljzJI4Q8LeKlb66C1AksJn3Q4y
2W+6MAE/SgRfzBiuvo0zg43CQwoPjM894h8EMdDsEjhnttM12+D0w8XDztWy7wmR8sTWpopkWOVN
jBndJos3Se842l+KEThB0xJpUweZfLDjFJYi3ErVybYkTbVIJU4cSWGL2LCRaOflE5B8WkUveLGu
/SK71ucrBVoaLmIQy8SZ70J3zxyGCTDFGFT9Zt4C5tgSFte5V790vzC3PYH8RKnHzI7IMyGpF10k
i9st9j7768cbqgRed2MslasjsaQIEfCpk/rrnxZpm1kXCIimU1dWZnMopNlhiKjBBMKod8nKQT4x
RTYNSbxs1CpMEBPLsi5KCHb16WzJJwlsiuqAytz2yW6PnJ0KNCBGVqTb7KL+3UBhj1RkVfk+Zwl7
fKZgWOz6mY1HYt5+G+Wsn5fWoZp/uUkb/GJ9IXMRrfQOZzVbaf7ddbSnB8ax5a1KdE6ThJOHo2iS
gn718Qvebqex7U11DhDIm41/Iy15+9NazETBz+x/LEO9fjLyNga2zPZVTbUBjgweZjz2lyYaXzUl
APvG25MMh2V/ocAHXRIefIA1PX0MyUS81bn80UvXfwozILNxZYQ1LK3ejnI17f6u5m62Z6ylABZ1
PCGY4uE7TAV6wkznuM/l5Rmpnwxzk9YSZSWS1f1IvFpnJJ0snk+i/yej0b0rFTV/ALjH309xsOV2
9Zu51ufiWEt+86py4cotBG+YXiF09JZYMJfGoMF/SXqAQLMngXRYRlhtPUfxWRqBGqm3Fpo0Z5VB
4QEm6XGqfWaOs2nEl5bHdFxWkmamNKz1rKudGKzU6hdi0ACdOyvfhDp3g2f3Rj1yhuqsFdXh3VMV
A4yo93n/LXpG/2uHUkZU2kf6F0gZaS9jbM9l2fbOzl2QYgckxKbH2JqZfBExZ7kJcA7Bz5Ei3jAa
6wr4Q52d4SAiyU5wmCYV2rgH6zDDAr9MRBfA+7dgFgi6D3QVGL2XSBUVL7qNylhBelSfMbe/HwbY
MU+sLGUhAKQZlbPutGmn9DHmLUy2h77z8YejvJ6K6BnILyoWgio1x+kVpxt3a2eOE916n06Lngif
/eEjIefv+3maqQxLEVFM20pA1OFIHdBap2rAiAjHWhm0YaHNEVEZgD22pP3/Ai6oq4m14zuItukp
EIaM5ry8qtGkRxU97uxoKEGLrC7Yjzv7MUstdcAec2rlUUWFIAObTAReXgKWqIhK4abEkOQsCy2L
1KXUe00O7Rp68OM4nJrA1o31IIHaJHbE3IVkMcx6H7i1p1pHfIn+Mz9Xx7+DpeRMfo+k/Anq5Yg4
hpcuNsrZotHrVFrf/FV2a0YmpkZ4WGu5JOzKrB7gxdlfCBkid667EIkNnvpJLmlot0uR4iEzcllM
WffwPSG7YrN/ubHNJvyBrsZy1O38n5xc7Gz528vMfkim5xXBteB4h/B4G58VbzF6JYz31wfF8o5k
sxHncdOuGnjirn8u7xAP8mMqcRp+Up0rp1CsYYHrDIo0o9XLPYKJNyNqPmOfW+1ogBVYTqzaZUlE
AnS3rNDkbyCwY9BzgPGtVYhcELt2pJufwIWQL6C+ZYYjFVFs10pnc09DrG170DYCKCIjNyDF5Qyc
e0yuWblRTIzvbTsj+sqMYx9bJL2sehnzKMzbckBBsH+vMSCgqcU9KVljB5cKGzMC+kmYe90klEEV
VOqZdaGnMSrvM1v6Dht7oxxB/PtPAGYgH3lWoMgisTJmXNoDWEzKhyOZgmBq4WSqscKAvuMm8ro8
Sdnv4024lVUD2UdVfEIzjoIDowMhkOxXSqqGaOQzZpp042/Y0nz7ejq5gijncfdKtao5J+X/9f4P
kRVPQ5bn5ecBDepOXUYb2GyMc9lw8mqotfu1fMuMvxuHP2ixv0SxSehHr79lKaJtQOGniQaqYK0N
datA0OgzkbDH+Ga5u61KDuolv1Z3IdhzJl90L/X+kN/zgAQ9Enun0VoTAjxAAHEoP2lUSzABwOEi
SfKVxivV0R4irr3tAn3C3juQ6ntEAb6lAnuV3lH+cPRKiJjDId7eHEgKx91DXyf+HU2anDArpuI7
mr0toqXatEHiYjqxOnGiWbx9ppeRj8V+D9V92Q9M+0nYzJt8N+342slyCnTNJJJLKWO2CVzxo8ci
yE4JlprvSuOlfEtzwun3n3jTA1bLzvC8iwwA9qKUq0ySnZAI0Zcep8h6clpMR7OVRRtTKdrx3Z4d
GghcrXZd+yow23BZhaU2SZO3vd0zp15HZhWizZqaGsib6VuP2o7qA+bO6O4FCSE1Fl6lOccMN1Jv
srkoQ6l7Nj+3VhNVUkrsH8EahjZNvgerq3ixZZDpqXzXi6ljzOY+xsIu/cbLKLCzqomR+fdjzgZh
yl6FRAo9kFolCwafC2Fc3qzJpPD5m7FOe5yveBC2ysII7Cye894yGuB+WQSzFYeuQn64dN1UyVJ1
BgxFflIZiVcgTqKeP1rwOgf1AXhyu/vJ02kSxv7RK55KrU806DLrCs8R1Q1alottDR421fVHw5Jy
MbAaop7pXnyD4CiU537NJ+nIlY1MUAc6cDN6oRmPaC6L5yePFI8DniiWKnHRDxfAySoYxfb1BkKf
IUlKlXLtT6XVbLekFTF09YvVsK4hGzMEzlG83hGHLPY8/R/W1MaweFxb43vT8qrx3R3F+tpQZa5O
Lpe6McAUwRGfCKCkWi8Y3+iuiRJ1UkQc2rEfbY7CEwG4ycJUh0IGyFaVZ3+jr2keAHoH+gOgAUXP
bQD0ZaMxLswAS1AKYpfryjtKpTBVoVTJ+Q8NWDwNvyUDzzZMwQPvMw8cR2XcaiiBcpe7Dr2+4UQj
88EazPqjvern8v2s5LnPaa639ma1nt7DFPN10x1sQeRafLk+fHfATsSNQn1TEmu5K4dx/qtA8YZg
FoXeZ5sKjdQIDOc7kfXn1K1x9z/Q1ghZmETk8Z/2HCTs3i3ZoutohXM2ESwbg8TBYNSdFLbom6rs
vv/KxpwFojIZhP1HjATENBkKCb/9YWH4nokq9Y7D1coxkNh1H5I4O8Fefh7Yvz/KPajRYvNqaXP0
w0/xa/OgIINAWYwrHMC4Cb/A0PSPd08Mw0ejU0hQvojz34N/aA2nSxo8+iISKQpyrKbs/k38z/ft
omSl2zfiIcHSJAQYjxhynndi/COhYcq5cGp//MuyMxhPzS5S03P3PrginKRUO+H8qbPIr8dUP0c2
bnb99jcX73WwezwXX9yZsVM4Yygz5t6xaaDRj/rBcrT6mPjplGWPlV9dn/IfZTqh/IIaQT58lz0M
ZL63dlmiWC6xsOvmwGUhJFHbrFC5YRwxgGxWnXuyBKd/IfOJaC4ePEgmjJ85DT79ntcXWo5rU9H9
VlBBKoPXiB7Qihamih/HnoP50Tzjn+8sEJA9NGnQn1heWKXMGwkSgqUE6mktX7xKLPiz+g72Qx5m
6edLji8ruKSB7ljdosSsijkn1DJJ3hiA7EKnUapCke78hXFY+Ymw1XfNppvEfmy3ukQh7cRYEj2h
+b7MA1508ZBudLqT2MkiRPFj/yy+nrBcYTh+92UYmPhbh37IxamCylYTivhb01XRzakj1nJQcfJ0
AMYoDEma7tDb1jjBp6mBwR9t2lVDFeWORfKpJPAEgfPXW/8n5VZy4MNUfeTCSuzogO6gQDpIL3m4
Mwm8DY57QUMZZDlFKlbeXDKlLIi+ciUMsNwNoKcwQ0HpVPK2wPGiLncqxgkyCcbtw6iJgLf7G4Lp
gZphQc1k7OQ4H+KbG+cYE3Dnn/l5mkhxizJwJJp3wpMjuSXOG4orNJQmBLVV539fpKy24uunOAAP
ynbrorFkoJcS1PDmWDAe4QjXS66OM1u4hjaNso9zjbCEM9hyGhe3ewoNWQWA8u3R4vnJWNuNKfP3
THhX9tO0Ms3kEo2C6ZYd0mfqoSON79ibGl8Dk/RI3TZ/A4vox/Ef8pqZ41fPtlhEXfXEmZax/u9h
qM4MUqttC0fLLQ3HUlOw3orxl8GN0ZWlU1pAzJxWNmtO+2+Lp2VxMOpp56rVEiMZ2PJUo2JSDKtN
u0MtdAPpGjlUjFTc9hsW0io5Xo8PxUx2F/WiJh9WOxKaJLhI8dzRfRJBk6vRX7fSWn5ZAu9tgnHD
L7YmfmiJfD/iNr48C9mDqcbHI88JmpQS9CVW2W9kRxFB1lfZoBaBxt3h/ym89vmeMHVp79/CmOaY
n1MmV4qd5m8vQJC+ZPEUrQzzK7tlgKBQsHcRSJ2oWhFYxZRQDZDeT7cyYrGp8ojzwjOWJJp5dIw7
ekJCzXkxBUZDdjIG3zsyWMJ1KUHknLHYd7giWeykN6eaTZ8I60Fvy4r2LsdLyxN7tB2R/1qsQ8uG
pUySoJCYxNeC7g98CB830AKwUBkxFZe3IfekLAxrvwW7TELBu7C1At3jUceEzTMZut/uXOk2oth8
WZSxpZjFdZAEBfRF7vTQaNZXNdii/Izj9Q7HjjiLlLNdIO9F5IrTMQ4UmHt/+8PxbeMCy4Tjz2GB
ylBL2vpfKhCxjzEgtmOQ8B8I/XBPs8dZJ2Set305PCvYRGFuJDqbN7QkCaYe3yHXcfleVF3Y+ZL9
qJ4z/FqSbLoTmco/t231feitqoBFcjTnZqTinlS0kMlVhbAoe7riwPJXsMovfJmYxqAFtH5WKwUa
GN4flYNF0mf7pcNA4691QcogrVdT88ZnvLRQxbEwAGtalTd18g73QTLX7cbv75CL66q1qIT8s+gU
LnAk9zq+egsdNYbwLW6VW0ZU9k3eTchTnuYW+QU5xv7fVD13hmqNDfbutNol4ojwqdxcH3eWFOdj
40oYVPknkSFOQk3d+XXrgwcuIb1VrNnHUMiKsxNjTbSAcwQOTT6QjvQKC0+tACfkc285nXX59s8U
+JJqolXDth/7oEgEgH3UmA/5rSElZphHlX5nFvRCfGXqDOLEE/CWKu/Lgvttni2RRmv7ohNPnZFo
zikPsUYMYNsGkN76MvAWfsVYhb7ZZZe3E6nqUrVBwOqoHhHTZT4k4WekWZ7xf8h2nBI1rGui0LJY
HsX/9qDyAYljPpx8nWmKOUvVviOhW+kdWdsDJ6OKS/l04onV+9lXGpmvmwkujTPhVOh4as35Wu17
loULVchYJtbqb79n4CcPWhKfbSNU8htheVJRlsIVD2o0kwBiw2TwkF+R1kSC/vHovlC6Hj8yWiyN
UDeUwrCBioZZDq/8hv0k4aLbd18pLhhqNNrMn5rbgYATnYT2/d25lNwd2+mikONdFP91fPbX/PvE
yXt1SCZ2ima6eRF7jT4KxURxEMpunsWpnCGLdy6m519KPEYSTAFnqUZC/YPt7r9daUpxK4RtfDhh
IzQYD9QxOgqdVUaZF1d/HiPgDJuDLdlZUxuPqLr1yGCmc1DorVM3R1C2zKXp64sHk4IMym6/pzTf
Q2UgdIXpEOl1viJLunnpXIsXjnwWl/F1+H1l4JvWI3B1BnhxaUwEOmviAdQX8jxj03ARSx/4QJsV
nafN2JnSPV3lpklvm8JnNFRCV/5QEgCrrlP2RX4XCJRZ23io0/UhMSJ2p9Tlce0G7ixeiX8O4gWm
mww9+3ohKgE1WBqurV8ds5x7tLZ0+gCBvI1+0nVr+1D4RRbaed6SUEEfBZpuBIlrXhsmPlLI9T6O
bsJD1Pe7iG16QIzXMEDWrVfDrgtSVtAwpYU2q9vpnADVXN9syF3CcizC1XpaKGRf/H9EenR6ca2c
A0gxBXKgg49CWAZFS75WRJWPGaTkyrqVPVFZWN9Wpn5o9Jrek7KM2VXO9tVVdOnynKSdnQvT+ZO9
7jClZ727S0x65Lu2tM5vhE0aici1MbyNwhs87VNWvXNVbRy4GRQybcEGA0/rgc+CKj6Mluw2B653
3hLGsTPKhbK1ScWvsx7tXhMyoaLRFPKR8cp1xq73yjY31jZbSrn5jb+6sWbkqIqu7ntA0iCUYxv1
akSnOFsRkkbs+/zlVar+Q3TVBCVgtglc5WoWWeqYomsJ92sQWqHNzGKaKLZiYTxwqMVaF1hN8kJ3
LBBmZGgoHzrcZhM/vRrInO3XBlo8u3V8nIJ/tHbSy+xypJ8d3eVmKd+wh3bYx3dcV+105Gk5vLyi
d9PJzPWJILXnWqbKMjLrDlgBiKMHOLbMODgwDqebse4zwnQkujg7/0blq/5IQqwV3o9GvndVhzha
/d5gcOJOXa0CPDjmRKTDTDAG5ggWlR+1kBxK5rR66swF+CdECud51HgyXmGYAYmtdWGi2UIQ/hCU
rYxZnnykt8jNv/ZWoAwdRRNe7SsmSGAdtdSZ+1QjTFx6yi3dylAAhmQsmmtIwQUxgkwAncJb1MTK
wkwsAt9/60N+QR5vfkzccPvY9GM5esC6WrcF+Yr4tlfqkLwyfQJNw8HdI7SWDQhyjVgnWpQlGG/T
1wjaMckgxPCD1wPZLwD9o4OaprA1hSTVbWhOOzzy1uGPgrEKKgFDzbZaPpFeq/GdptKfoDcK0q9H
RSzICOmhjaX6ehMklzkrxAGn/G0/3X73Mvyrfz9ofzu+aNBrJO1ymzErH9YVDQiK0MTwMQUxEIgb
G8LwAmw2chd/diHzF1pxaUniX518f+5NocOinRFYih6sH6SXUE+TqDnBE+WM53426cL/z2/3PHdw
PtUU77myJjQG+gjU5yRyOlrbpYPeaRJ6t7IGgDccNyjla/qjbeMx2Tr1WnzJGxc/3kfYKglacqT/
WCKNDwGnSYGVz/l7jQ2W9DMTGWbxyXUpL3dMo8NXLrHh25Buf1xWZB+OH07DZ4UCVrJ9Iy6Oct/j
lbuQDYueRuAiTfieqy48PppiUee+CFCOLqyDas1vyOwqpanWFpLy6ulsm2I0LS5DGmlVazdvlZeX
DwKSdxlGYAWDDWRkVK5xkdAErIyr1OTx9Viaj/yGh7RTf+ko9C2X1L5+VwL6WrnfuRxq+MDTjeh5
UOAmvjQzMbZ/gz9vJQJMTfrdE3TavGLdVZ/aWR7oTp0y1V8QGObZZnio2Fnaz85/SExFreWmb+/1
w6Q8jwGTwu6NVPJm/UzhNR9yCPo4edyXSkN1PVv7wTdPEK2VHTFTdxmXMFt9PrFBhY3ueKkYoxo5
5Fbup+eYuU9o4f1Aw/vCHeoZgj2UXXqydXoe2V1tNZzD+XSn8EQIrMxDnDeplH3QOgqwkkhR/ae3
7gNtavp9A+r+ZYiWhgXIoHSfDlC0lheAUvgtVpVM+Jk8XhBQL22VgJ27ZPEVoK27hj5jcjctpXSS
CMPgJ40b4k82f9BGqXKo0UP9oXj8nmX2c28X6CB7gy16yz6WaqeWv81JCVGDO+xrNtVfnEV2DZTz
HOEDxFdUwU75GT1AW/poZOKjZDwb0hoTWwLklvoAOYBoed+0cuN6ZOHn97xvUKUA98CxzSCnGWHL
VcOG8tfP6kYOlBKTCKX7JZdMIFoTrJoUNmf6fdVVQjTPCPdIdHdcOYgNIG2+/dg47h/eaQhcbbBM
JThQSiUlgBFVWVJh/kA1coPFdoK/ICDJOKDipd8eWIG4VSd29zI21ORq3zPXy+AIalLixTt058tj
FWam97BV2XC5ENL7KsdsymW4EWu6eXHrsGcWUwOhNQ392a7cpJt7DxqLqsiXOXK3+ZnLnfckqWle
NxOmb2pHWRkOZQ/zWnnlCqB88ke8SMHGO9OCcjUgPfpawU+asUP7chGNiYimYgDMbZ53KazNwbpo
t0FmUKT2uw3AGzxYZqquhp8so2rJoRVhBlrp8QRIrGQpYlJmSJN6SLmqghgGqir8TGYbV/LV0OS3
epc9gms//1Xncz6aOVshPw9ZWoeFKWRaEJtO/ezKMx8ZiULxtHSMFkizcY4j20gMkt5Q4dfLcHmE
3Kv3/WX8ECVtokpn1GQZmFeUheFwKzoY8UxZtQBCNhTeDjGqUGbllqb5qhd55XR0b+Yd30enffPp
DC68W8P+riWU9OJ+ITdlvXGvlyLrBGNb7BlR0YQKK+ih4txRNo+hzpZJHlUvMXQsHw2Q1uxrQuwJ
pgHhnYHuh3W0lCaDXgnWzi++aBbXkPwQ7jQPy+9y4e2eLSl4evbrmcuPtB4vNdmSyPN+Qdbsugj2
Xcy66G+nAX0ngcNtXL8EvUK1A4SkNndVrxA+zvr76OQG7euuZWRNOKaSK+BYlWAeytejFx4MVRqF
m18MZv4DtsbLu0cNGPvI9XICTR/UlcIhLx593cXd/vUb1aB+QZA06ABBei7TYqZ2URtQZ6fZgWF6
a8Kt5T5eueEPHIfFWrvABydSx3haF4CZVC9z4q+dSiUeV3fKP+35XIIx8GYzVbBy564UEV2Zw/Gf
c0YrwYgPuREUNHLqndBVioOaRqEbbF3OJYz8hUl9RXuky5IWCdi7+FK1Ip+Vo7EG+r9qx83XhrpZ
76ws2gbzM2n6zDQffN5WKOCQLdmcJM2UK5z9k+nHSt+H3FH2P/r/22NhL/9dx6X1XxTtPzbHTwZS
bRJ/1cZ9LE7Msn6GAsV85CKGCYMJzolFlMHrz8AnVe1kIPrMBEHBOvG1znvY1DzsQcLodNv5l9L6
OKJOKQ64HFZfStQhDnLvk95rH1p+J5xiOUs8KdX3BXW4IbhK7zjhHhizSDbPqrprMwXJynLzm7eI
t6v2YLNk7sOA1ujbx+H6TOeyO0oGAL4UdBHijp0hjYyWuUKrmbLrXCvGQprjWXPc8/YmjOmGzzsa
1Y1E2k+H9P/F5zfYASrC6PXdj9ooW2kJPLF2liTsK3NP1MIhFVNthozq+1oAUjtinB9PDd0R1BpQ
XAHdCk1+n8QhpE9pKHM8mfYD7cL254bLPExMgQtqMYcl1GJfklfJf7ajSI09w+YRg8mLWqRpdU2z
f6pSfYk86LWVs17G/iU3aVqM+ZYxcLwM1GASRrIniC+4g5NjyWtaIICJD0k9L3UmfiHQ1SsRcyc8
j2Dpa+HaSu82BtzMVkknj9CNDfHBmavNXqsN/vQtKA9sTSVQZwDM/IEN0v1rZ9uC0VGTdlDzT+sJ
adCKenydm9AegfHz/ELdyDmVTVfVvjpR8aCkGdkW2Q3BlQVuUMg7J6MnHszgMbTJItFsTH0bLhju
iAdobLizQS2GIXZmkQOfeqcXKdhEnPpxJnRaLwISxZMeqVrqSU1zY2wPi5uidkVlEKpKGPVoxE5k
ur07qy/xGOrj0gkzcK04Fq6IuBbBV3M5qGfdhwzpm4voQWqDFPnW1NftOMdVOsuS632Ih3PjlU62
wwPsU4QMkX1W8rGkL7rRnWUTHnMi7wreUFj7RFIRcQbmtN+USljravYid+/L21jA/AyQicExkPgZ
ROWJYyzuClpv4AOXPpzigXSTmyM+2TxDcvFSntFx6hT/drXouEuOC7nHI8l83qjfsNdJ8+vBhmSr
kRwBhhfnWY6iZz7DhUXJIN8Bzb71JXEPvdYk5rMdJTD86UEwHianfCIwan3eICrTMlPJ3ko9RqAR
0jMDMZZPm3LmDWzySXkVGpVX0jH5QGV7EjHURWQWNzFe+4pPTdHLgC6idfTEaGWv3eBbZTfpFcrB
3YcPRK7WK29Sgx0JNTKVNIyhUZ6Q6PfnjFLdwt65Ruds81QZnGx1g+N7UuGQNgAkaWqCpyNdy2po
fQo6/NpHeUTivapeSRsLDuHWeZLpH5XMNwoLfE/ubtGucJg4uponfBOrlcUISCqKFYxjpwC8PbrS
ubF9vRgyTniVF78a5Kl6XjHcY1xD4Jz7RfZ7OICpscnZACEt4Z5M4cGTCtT3wuCM8Ac54YfXfvtR
SsS6wDBLX3dNhH2BwKi4A6dqtGRJwB7KquhBCsS3/SFW5KT+2/QfywFkMKe+2NREkt5OZnFNCXuS
zxQf9Dgd/dxNgds4gNmZPQXRhgUoewHXKqLv/64GM5onKZh4yUKyhpEkunhZT7hHVWiZZzKKg3us
LAbhd8dqMjD+QaoKOx6cacmj1sN4F9Z0MVhJRdPT8U7cTqUTyvRkxq94hKfm5EJnb5lldTRWB2Dj
ROCDfAR5d6boD6C6qE8+3NwrAwP1CoQF0TjZ5gjWZqJcTCRmWUqPNkAuyvG3LZsu57dEi329OHqw
MQvCjTU4J3wrw8MvUXmWUf7Mavj1+EphCKxD438ePaR4N2EUqa/kmlLXtuJ8SC0tSMwr10rcPQt8
cQs6Otz63Hfw30yuHKjh6pstj2OolKLYtPTzL6iBOAkYmrTjQJegLdB8gWcIEKx1Bcmstbuo3ZDB
PYT560wT4xACzakvHH4CocJhJ+mcbB8r+pxXBiXj6GViufHhDyL3CKm1RGO5TVHX1EBD2IuLSKeI
l7jTf2RjmuPQmm4NyNFVxGvkWOXXIzCYWHUX+YW+Qj2QTWrgWqP6SnE64UkH2mW/wgpaBR4zEtGi
yJOmM5fqYws8OGiFg+uRNrutc5nPQghBV89e2kpTuMfYAo8JFx8HYq6xxC1xR3ZCMFdK6n7z/4bD
oJrnd8zBa6GHsglgJlPJ1ihPe9Uuktr2K7AOdAIWAXdlu1C5QdXjH18nZAkEM9MtdrxSi5q+UNWA
mYWMYOkvFDl2U5FLUoO/jYTBIMtJ3/Mj50PLg+e8NLm9a5s2g68+WJ9O+hHmPvToj37mgluXScqJ
hSz/wx+6dV9TivuRO1u6/rkjWHB4kFt5ZMR6m6kkXwUIN9rOX2O8M1XBPjnDmkWkg2xyh10mPsTN
3QkYQKXisb+KkcnpHEycvY7KLKu+Wfn48N6gC5vfJBXhbs0b/P8yxhO8oFDytH7Sd3AqodWlS3SE
ZPFVjmhl87C1S0o+kz2CTWdnqjMgmmVZp+5dRgd7rzgTZjZmM1Cqdv9mJB8/P9i32+bp9jbxkYuW
oZz4DXnlg67coL8JtGuaQpGqiHvn9RUolY09LWuwdrgEQujMexepNlwowBCKtmpwySSfzInQwydh
xSgXc40PY5XVY4Q715jfc4lkVmQ4RCKKg0NPdwVHaoOVC5coOaW5EAXuWwb72/E+WO9x5d8V5FTt
FCCoORoiCBhiOMUYnhiE9dzlo9+EOhIe9bqgvSVs3IPj/0XcrvqUrGKtp9Q3XLx7r6cmEb4X093l
nsUTuydWAtA28uNtKwg8QpPS2M8itWBxuOVRkfO13HzoJwbVIrd+mwcQMKjB8n/1N8fl6Bae1zH1
d6XMuZDDFaTZHozlJ5qrTDHYPaAu0cxGW5lnrczfAEGVFn/Bh1QkDYZkjb6Oub8R5fXHGPsIhz34
cZL9I9CBk5qWgPx3RahH8gD/roXVRhFAFQOY3lo69PohP2v2yqujYstpAxk4vuLkb6iBi8wal1TN
Bg70ScMmPQ3In/eG0UESJpdOJL0zHZ0kFF26/HJfMG4q2N7wGke9nUUVD29htzmyqXXE+9mlf7rF
2xVfQDwJa9JDuVQxU99gBKqbt3y4z7/0or9aNXqGa+T9WTpbShPTrz/RdU8Thauuj7RG43n41gC8
v/vykv6EGkcPVYFVj7jpXhK7zR//VhBxwQFEUoi3DkFMQjGeRVnZgU2tw/ym0COKSVS3rIjUCeI1
IbE7nl5iyqR1P0lPQvDH6/SlzoYLFSqciXX8QvgMPHaFlMYhfNPv3BegMjHAXx8h+674SR64rMQ2
b8Sc34IFKrC6fQagmWhZHLKJ4wOQzddSw6zVXiYJZ22YuVp2B3yedkSxsbP+dYxazskO1kqDX/5y
dbf7TkAZ6Rzr1V2GAxpkgZvm4lAa+zNT+D5Xd4T/8uZfnusbadSg3fyivgidTi4s4Ij6wS3LbcZc
D0TGKuXAIopXrg/pC6q8dd2UYkBLpAWfi3uGUwh4JOcj2Tu/lLhb5rYaE1ovoCpZQl9dLWe3WuE/
dFEQTQUZEsQWknhceIlI1U9x1puCXCznvo2bg0CZsslzP/z3ZlWO5Ye63aMfUlCzBu3alzsMPMrT
Mm8zTfs3CKYrqGHSbhCaUWTIL5XrEudB+lY259FP4Vej6/7pSuPNEQqbxzUG0PjF8QLjIcGS11nx
xj8gjpmHdubZ6/JsypOg/SttuSU7VhVmzyl+6QRMZW3tatiTUrtx6IpGwnw9e9lAY88TG+ssNoMD
q6zeKAkTG5zlhoY/hy4QfI4DXo2sXBixfr/htgrO5sMEMwmc5+/MTC4N5ouZLHAnnKqa5jwuhWGF
GS3t+gsL1sfGIGGhwUpClAgBEPoKCaIPJegpPkwDcIXl+sPQFL2NxhI6XD1lmGsyxfXkeI2+Uw6i
HnSwmXO0GORKxnIGkDMEYX+Kck9YTFRsdEUgPwIaqBcW+OsKmTjzJz7IivgaEUUQF4T6ka4MucVu
VG0V7IvckxZd1jzvGzRKiITDIFxUHF1bvulB1OdjQt2VyodJfQyYUWDoVPbgj/RxDR53uSAjeZ1O
AsKvzFpWxWfokgCdrYlRHA+7ykF7Qi8TzakkdwGhNLgt92ejNr4qUdrqHqDAsK8J/W5Y3bhdANNz
MB6IIHZKaDhkbMCFW9RokHY2mBZghMjv+3t61nC61o5z+Z9K4+D1OOR0r3/dmE91/v/g1hkNtwx/
rZ8zZMDGjJjgpn26Y5J99O5DmAQetWVTlPz5d7D9gU/vLA5tmush3p9wnggK+c1PZ4asdSS+Ar3S
jVqwlQccFVxtt4kAtCXVda/XkD49QD/EidRLtpkhgtlD46ZWyQeQyv1OlS8eNNtq7lg3k/EQHdKH
K6i8roXI0kVP9XIlM4AeUjY4h0wHr7Hmexzu2ee9CGSfngrQKM7CSHkw5Ks94dK/WI37dOjnU4U0
l46o0ZBv38aNZa3NjWo7yIbBIsVVDiQwmFGan7zj1FqoIrITX54piX8X2HK4TUpLeuHelIjvCLGJ
zCVoZiaNt0zOe17ZLgRYUmLWe+fGNE8Dc6kiCb0akgnpgCgHooQ7fPygTt8yhi8Tvex5llKWARyp
UJGAKjfThix1LRF4Y4CYMZe8DgJV+lo0RGcRQDWlJBkbSmjVH5c0ucT2CVU0019RcouNscjF4y1B
8Eb+m7M9l/w1hil/Nx2UlchM9bn8C/tHjvAagOHGyJwsO4I7FPXAZhqkeaGuZ6CBgRM3KIIARCL3
tHAovxkmSRBqIkrFSb37s4McBHdT1WqNq4g7V+R4G/0BlxddnQo5Sna45EkmeJTDkIYgN/6f4TND
zLngydBJ1zehEoFI4AGhNYaMdLkD/zBjCRChqbT4XIwnQraK3z/gof5pK3rZ+b9psIdMzOlGJryU
5iYU2xAFksjm+4coqDPdiToOOpyVXNVTrIB2fJ17r8ExN/wbB+ePKEpt2kfF4l42EW18xyAQr7OM
apxEuKVXtI1u8duJ4Z6UwpfLIJcaB4xwsT/LIWmfOV+b25hyikTBaUI1GQvveXDsi2PktJ4bqZG6
w+oCKF1m1e3Gg6s3AOwRq6v1Y4x7/lMLiQ6qpDM3+HYpLNTOD8Im29Tkwbsm7oURGI5ykiM0kgYJ
LHT7TbIzM0/BTLyF4Y6zVU7dEIgtLSSW+d1xsMmCxXcX3d7hMFAPFKfHADPWvlzgQiLk1ouLAkXe
d8xvg0jYRCihnD6pjpNVdaUQLz30DdAQLfIBtF0VmzVesaSaxb3xWgIPGmsU6XUUnNmvpxDcKHVe
Kq+kc5aH/Puya95dU/+HLdzm7N/FGIH5EqdZ9rspkoHM7Q1QYZVx3vTT4wi7G3ZLIEI7yg5qHa1z
qpJtwb1l5QMeUU+jXBLTjNV5OI+3FQpYEE3A05jfCWN36UInv/7P/cSf3OIQjx1BKhI7sewrQ4fh
RvjjMRFDIqsN+OlFYOE1jZ48uwFf1r5dVP6NJ6aqJdC4dFxtBj399UKZoV2pi9hsNqVPHfRntehb
4D+QEU/lXZy0cyuo6b8qEl9T1Y6lzt50z7J3OocVm0AD0WKpNXjtI0LSwnIEvthdGoB9FhNgqSGQ
T2Je3meNLl6AoRTnyVMUTfU7ycgBZ2wbXpBhedYWV21J3Y4WTinoxe3Gj619LQJVkcRnvs0nkUy7
3839YdokpNpIlvP8MC1MDbhBF6+kLdFCPmD9LfpYMzvPZH4k0D/rTQv7X5Q/HQ0OGTu6jmA03S//
BTG28krtJ9SDKfBhH+IdvgN0wVBRT0MtJqq5OiQsaW3B2bf89KfiVarapWs9750sgVsnf7Z8caoC
4eVyrw7k0scSH/j9pGjfJF4GEZUc0sNVRq3tvuLbKx3CQSAVwfulKi893uhtWA2mSHQcwd5T5wgT
cHam00CEW+yqOwWF35z526JCA8OCKeiWLp1Cl46HZbZbEklIk1RSzhffbpDHUO7L6SSz5luw10pI
u3UOwQU1FiUNvWgn5oIkfz28vYD35xttD7o0T0wcke14ojX+tLlCUUtlGDuINicUDTL3PYi0Z/ce
RWamEkK8MznArOgX+5h80Gg1gZw6cIzLMS2/8LU3PMnljUtIspX+vjSVbEtBpw0VRcZplp33Khy6
ynH9Ro/H+F9+Fg5UkWzOqNixCiLIZozMdxJRt0TqLWVm/9MVpPb7CeIeJlZP9ceY+Xz+NfdS8eJV
NvqzH5F50/skEennWrro9vCaotnuUbsLAacUMxjP3cLDFLUQHFoqmwSuhJQjjhiX4vFjp4/pStCE
zg28A3THPo7/nFK5xCLAbRRr3+5y0EWAJw4SA/NrbW9GAX+texhpXrD0SOUUW3NbiVYlpPGlLeRE
f6Rs5DuR42HR6O47O8VIORVaVbuEbZ1i8wte/0Y2gVZS/q5OqkY+unF7Wq+CACd4DuMp8J85a3BL
CPOW4dCx+u5WVtU7eC50Y5VRMwwEAHrAcCNexSUWZyxcoWas5AlVkYWHPMryZ5i6dVFPJA0nQesq
LQkEKUSVlyU1HcKIWsfVQeoMIiFIYY7TIMDHS0Hy4upwBMwURVakFJPCmUxLHNWqpsU5XoGkQxaC
N/90VRXRiapwyxY6c0NY5mT5VfUCfXdbYYrt5feXT6hokxifHE4Ua074If6vp6zQq+Wr4PyY9Xab
lcI29FPre7oASEMEeZJJX6UuRzokURQQRDPZB/aseSTjjbhXePXLWNEExVvPKhQlNuhVJJv4LXyn
4Vh/mXSEvomYbcbp2aVQ8CvaGKEIPwsih7rC090hdYEWo/hUxzrmXnah9FD7Fo6E0llzz0uXnj8O
gC/v9AAuTAHdWOz0iRw/rYUTBIdB61PkSukzI+uKhc5TbEn+iiI1bkBkWY90w7iQo3Ve4pavsw//
uec9gaZyDJR4gVtIVQoBsvW4sDq/103plE6WlB8zhn6fgwXi1jaCCQt1gL/RAjP5VEMXS6o48fj3
IXbQnB1uzp4xTIsPaO48XSfkYCeKMIvrS0tPXK4+85zu+DnFmq3rQpY4zjd9aFr+3grBqw0q4f+F
ilnRULM4N3BoyLdt5bMDtpNoicyQhr6w4L9SwvHANyaGsrQdBg/WoYZtky1/HgkynbVter3OKoml
ZvqmZffNc4TNtuCgBIfIpso+sa3YJvL1SX3AHWgAHRiblqS3/L4HRNafP6IO3r3aqd8qJA6uQb/m
ct9de0LBOIyIfF9PB2Rv32TbFXmb+rGq1Diy/mOn6gO1Z/JAaGtxvLq0BgqEIFHPumVhYXP9yyHz
ZSJR613Fs6n+lFSmYDFDlXyjl4EAeAsZH8URMtTQN+ZvzRhEZFY8fM3rntDn0ETUx9RnA04DyE6w
DAE8r/sWKitMmw7VKaNx0c1RxJei1ZnthiEU5pejt7G64PYY8CCvra5AX+EjtnvRZiaBPG4bURXQ
HhQthOddQALDRDR1YdWAI8EFY6RfU1wMyKNh00EmIBRDFEJa/m8N3qxRSekp8nAcc6dY+FGfmsP7
79mK843yAWfIlX0TChQqbASMqAeej5V7SzhiEVBZMTThQ6ow0a+7yDZFtss9Y/ppwYQeCbFYAeAi
0AyoqR9P+rZQwarhEkyvbk1uqyuqst/uak/3RFRDKDpgh01Uy3IoEOAKf4GU/0cSyHw8xrhDvmRC
FQBvwkvR9lq1xdMOa+03g8dP+KYvDbseaVcXz5+wZNeM0M9litBuPSj8WTo6Ev3wW1FthVYnIQ6l
LEFN2KVKDNchemOTu8omomm1kvyV7MP07eRI1xOicZINZoNVonkOW+RhPI8if1LMBrqCnk/Dz9gN
w73ffKN557ADW4cHztXdOcEZzFlWp2AwIvVmPcbPX2bYaMHhmyUNH/eSr+dO4vWaBE34eBPZZB9r
T3Jmkn7lkROXtmzpK5qt84BwRnUH6VRKIpqtrHjrmF9imdouHLVyMjFh/XoAvapX3auE9p440B9V
zLLYinIaf/f7FPJX4r3R3so9bp1qTVaPbvMRqWIp6cVtWqMSwDh0XzPQvwe02U7xQaI1LYlwxnEw
1BAXy4CcUuEev4AD0UswD1vOXmGaolXDt+SihQsYQyNRVBXZ0VbLt8PWKS6OAfcrQ8o05s+xH1U5
nkNYmL8EpHReBw3RMgTplGiRNpGxRfTvj2ahu5u4poliMpJcVcX5vWleZO8jT9K28nBoSStIMplI
ipK6m8ROxTema9jgH3Poaj80qfAuW2ojJBHHCNQtoRdbbYf+w3I0sGzMev/P9pSBWT6gEpB8SdbU
qY3My2XPFWOgCwsxgx48d+zaHa/Xt1Gma0pKEYbOrvOEaI/QzqPVozrwIFFfO75n9prz7El1j1uF
Iag2cWaZmu8sQl40NdPgIUNOYrvA8DDeL3R9LxgGHKyE2atBmMH6gbryi+dQz/2yO5O7hFbbEhGU
T197lomqAsxp0giqZvTu6u+EKA/5S4WS67mQkt6RqwowDgDmFtbTuxMQugjSdMQ00LIUmSHeHJup
Wtu6Y+JJxLcnVUYOnIcAwZwmiy9h7BzGiYvtsqpWEtyFDGYFHTl1dOZDQuHTb5UrS+KyEEsguzz8
Dk6dOrRkowkXum4uqQ7tlCctGQvI8FEEmHj2zi7Cjsv0b54NbRuJyjwlhH8Cc63nYaUvVJ1YjW7m
oE6l1NVuKU+rFCmBBrXdlgyK49eWETPtwX0s4cQ9JIf9GL/GosVV3STc6KtvKu1IHG/8uYA9D7AV
yMzhp3skKWpiJhndyu8RGi72bfmYHVLdZ13BfHyuH7Zd/HW/gmWP5kb1pZ6uu99dzg4gcD25bXqB
VwyzUnQ+zNUnyVlJAq9rH5MCqjU2WemwrHsA/DGLudAX/7wNDiXPO+Y8rSkC2vJXjxChIm/FtX6H
MOg77ftjeudNldYuC2g9XddtY80yJ400cYw5Cvoi0MIgBwGCKpMj/wPF30Z8ZB3+bNpKxApqVcYk
UtELMdQRUlnqTkbB/ZYbaA66rOHVW98EslZ6OP10Swx6Vce40jvlpvnaaJDH4IBgktDrCyhu6Aue
5DLrjzIYEZWZtlR069HYGMT+f7Bmu6m31gKAeK+TDE1kC/GUcpbbxRYg2AdAzIkLgJiY9oeJCQtn
9h8Vr58dfbV7nTgUpiyxbQr/Fu/zXymlHWJRNYRTjODnVfzdIhkXApDzqOOI6ks97oF7QYouJxAB
A5DfRNFbUkOFomYM3+NeZTG+7NpPIUWZ0Y2Z9lFnQdKWAaPNyxGez7Z/nN2ukYl5OSVEHPlPBSWA
WqYEV9aPS8mdT9kvb1ZMo0xcLrPLDmhrCvFYjA78pLAwek3wf58Vnw/yIW17Y/KqgJUYbvxUqW6r
7gY4n6vdPAlIl2Hzqpexh3MW6mRnPF5UjfnPlegWLVX1SkKH1JV+Zf3KbWCN8xhuf4gYupE4aLYl
Wx3DCdQl6+3eywg24T8Io0Zqa/d9h3oZhP9rfTzAUpS+GYdfEIalBWQREPl8t0xuxsbqpWh5zxHa
AUHR7f6wIxyaYRTlOldX2Z8SPciGe2Z9QzH2QG+mof+7rH8n8piUIQkW7TMVAjrEuNZOpaKMEw1Z
XkzjSQrqI+5j4Lxqpm0ppQ6IupeMj3gem6R9qLZMXJ5QmiQH0DLcHBZWaXwNVlmWsgAjiJMgwhRb
seAh0M8nZpaVyv5PrtOS5H64uZZDdpPUrqVnWsz+C4inHk1ow7PzGddfz6Im5WZGRGNJsiU3uw35
zulPnHknJO0IoaCtvO4wPp+G7/G5j4ooVX1GhSZEi5BQzmyXEOS7bxVabMbLMjdjyFElOEOqXG0P
cJ0ECjzMZE96yQYq5+2LuFfmvm82wZO/+1J3VmisKQB1SFqH9Sj9sSxiQGSXS3xE2xwsOWnAPxHH
DBsDk7ebjP/wlyO9jjNzHdd8D0k8IX4OQ630E8V71LDKKykuzwkTWJHZrpUE3esbT5g3/0dGYDZy
/TymdwmH0J2Nu7kEF9Y+sTYrkJC0HWANCwxEnjkNuaGwBop6ZoJs+p4xJ7vcOTbemeuwVoXEsUuL
UsJ3puhroQd3h1BF5igksXt5h05+R/RQOpBbgnAR4vQFAKAVhnY+Tyk1kPSSabYp3QaX9njUIoSx
4KR1tqWl3pRJSUUQRKdZG3rvK7gxtZNpPTT/v+TOtffiHUCafREFkIg87Z0konnKZlLMWzBjIorQ
2cUjDfvLguomUWb3Xv0NPYq4b6xB0VV536SagC0lGYd0lWQakMGKA/3XutP9iT69HXW6I1sNCAST
cFlcGTaop/OqstLBxCdcK0XFfmUDOUp3uvrGudIOSKiqpCjbAZJAF0riniO6q9ztexoJnKxp+krX
WGOI5ZeM/OwaYYS5pS8jx0MCvA/1bZtE7xYXwzp89gY6ArXAvuOWErEhYF3klc2MrgRDh0rGC+QO
2OZ3RujCKGa97F/vUVy2F36k2/x1xshr/4W6VC1BuS+TEJQ1kEtiy0dbB6DSiI+/gvxb994nTkfh
O8FlFGBDP005uZHDQLW4bwFP/Mf8P7/Bp+Z0MUiR7iHdwNelMvc7GJF4u4hbgcfXTYNlspECEP6L
ovAQ5G6fzkr7KpAVbE8gqQqnyd6yUem6wRCTAM6SGWUBW/lq/yXnalJALrVJbE6dIIAGECIjC/Dw
Uoh4dXbkDcSPR3dg19tyWz/AAK/l9E2Qig8A1IJxPmbJkuyJykMlD5yDicAhMdSaUjQVLBkf0qdB
mUkK3uq0yWfgDP5QbkRTEsvSNfoN4v3BQq0a0Yvu7xkiDrC8fGNhdQXho6RCdOWCXLEn8fVeUoNR
wGeeK1ZE4LnfErEymuFke3E5DbpyLbdtTTs4QQotX1sOm1qnO2bKE/jRTnH8CHTal88LBjbjAZsA
Y3sRcZt7zG9XH/hZvaX+wrk7MAl6uBRDbzygW+LjG5gBVhTbZAKCuXWcsVtpKYk+sflMa4vzzFo/
bUI+sX0DkmlVsi009i9OILyoDAQcdqS9HYRzuIvfM8OlDKnuL3/R+/z1WRqJres/9Or3iMi0/Ozx
E++KrviWsD4Di9tEHte6zhKGyKTeAD33MWBph9KXqS1eQs1x/vtDXivzvKbQbCkPjGvvFIUemm1M
RfGSDbF4RSFmAZcDGcjdpub+gz0mtmSP3/mNXTPdqATlfHqKjtU//Lzlgq5MAjvF8MBeMJCUWFjZ
st5d5EP9rFtDykUU83v0NIfSqiUSI9W2V+HALCEKsH310BawBcMwTvrIIwjXPSYBiF9Nx6iNA0I/
ZJN5Gf9vlMw3MIHiPgVTqtSJ6HPhNHrK0XX7oL/qIYal1HBzTdR7/TpRWaZvyT1zeZBmY6wX4NnU
W6DPTq8S94AybIl1cNr/WcA1z4+vF23gYtJ7oKBuEcbFlxidFFrvouPACkF/psUjQ1wQ+7WLgvDn
3WlBFtU2LsabQVxj393H3knvRIX29a4Eh7EIuyOr+ia367/mL/VIJO8Xmd6d7fPQ77SCpEJWweUf
i5MTI+LdniHBDSkN/mbhhS9PsFuIQNfezOL9QqHkgGFS6jZAC6KaIJqcmYCstQQZ2NZGJkg5Rf5a
3CNECJzvJXdQt3bmdiG+UMkqeKCcafG3CaVn/eg0SsXC8PXgrSkE2LcCq+h/dxJxt07W+5g8guBC
08kf1Z1we69kO6ETUkE5v9Vikv45X1FQJFNEOu0h1ARzXljgOpnHPFim61C5njV4fHdt9KL8cYfP
rE8cqWNDXmbvatPBSpr3hMVVN849+A+xHD1rkD/6rbwntcLQPJZMRWPBNVXuY4Hpi+8VAmLme3+N
QWFp9QKK0HngnE8oO7HR2PkXY7vgSUFZXaJg8YXE6cW9bChE6N6qokSZpBV72KAUQXHQla4mNM5B
yt9kdflWTKzM+QJr6Wpv8QL/TB6i/92gf3ceT7l9oCC2ms8VMA3p3slYI8aQfzxgawXrhSh1yiOC
UdQjMcZ8vBvHvKnQhG0kDCUUCn4+yqlud7ROiDon8eX5tjQKNo4IHXNg92hnKU8Oa78rQsUuPn94
kp6ob/xx0hH0iASxsNAIjYLkgqEc2hEubv0hrJePa8RRdFXWU6whSAYnUTITkvhc8H1yNzZWsBjo
r24S1Zd3vQyTtpT0r5N/G9IIC+vJ97ElcpyghX4okOd+Skxqfa9frM0x7RdgRJ1NkCC48QpzhXeO
Ne5WFMmycMkpZd5iy54mfgpdY14AZaqj60TRJcOWJZ8hZezBNs4TkX2kRODhUFI4fO+cZ1BWtW3o
hQpWkwIBBDblVSNRe+8IKVJy5NCKkwBdxT8UhnFPCc6Rq4RBrRSpoYKQBqxLC9SF1BH0/h7YMfdc
89B72gQ4awdArTpYCG5MNr71MUSPJOG5BCGeYOtGj9mPbo0B6qkCCug/p76yycbPq8gnqqvjMAdZ
a2oREjEpb22fgMALIl5e/wuZ+xKJe3zvEVd7sCCT7OKmMVjyWVFDLucUWxVjoQWiAoBNJCz4QSWU
1SiX5L58BK9PeRATRitEvJQlJpq8Tl+KJ4VXzZq3tBoCHBb3DJrK6PW8PwB8K8zkfW4Cyzxblbyu
kqc1oXV2V/JMmiSY+SukZoJrF7FKbNAA5lfizN4Ns+Vo92B9tKQZLNb8cB5TqTFxMqRxpSJSC5Gj
iLOJFVMjOM5Cnlx087b5VClvphgnGJyRl+q9WfCBzVKJLeVwHXrLpY5hBkRWm8styW5gpy3g+1Ct
dPCCxb86juppooE85sLhFPKLbfXx+iRHemFSNB+Ihlk2lEJaauRnR87itafktUsnfLTTj4GfwtYt
Mw/feZnoF6FCm72sEFsC5iY9YbMJe3PXDF826lkfrk5zy6Wwp5uDscSGIRBWhPVrkQ6wDrezbJoB
sG6vpJpI1R7k0HPA4XMx1wybS6+4HALD3Z19WnO3N3OigXZJAEOv4mX8Y3aciwqVkw+yKJXzi2Zw
RYW8L+o3eRr0Bou3C4i5pHDxf2sWYmQdotSVswKBQouPQyjlGjtiD6LguqiggZUbC4DXUyhuTB2i
ef3BSyzIoQmPBUE+aDR9wncOn/M+BViRmslL/1iSRnntKJMX0DXrGsmFGX6+dvvS+RdNRNAbKYgx
C7hrftEkqubeOsfS4ezmnVAo8D3cGUu7Pj06u3tcNjXuEmuteARpBJHXbdRKhiifkaI9SRaXszO3
hA9hVPBEuO3E07P9okCAJ2haWqveC0hUVAtSg7z3hef05J8KMgt6jpqIbsLRJR+VEXyodzNMrWUV
fWbGy8OZGM48DCV1pd3VoqVmrQzs9VsE8VRx2OWMAaR+49Vp0Gut7OjQTJ8lDBqNIY09Boyojdhp
kaOwiDwmXsyqjdP2BnmuRKj69hPo0k+9WJUCxyd0MRZ0eN8yMt+I3h1aF3phqJguEUil/NfQq0Q5
Ubgjo2Ext6cw5gmq6iMFyzs575wythpFcVKCKKSyfrgSFLbJYy7KNZfiTXoyoFuu3CG7acjh/Rsc
a3lhKsfRkTeap8znHxIke59wrhDAzCyzHA095GABFOtZS/vcJevcde7Hnu6N6PofIBVnJ8dBrx8r
h4bvKWI8evqD/Oz/L+BJNjbPr801sDUFpvcfxn/M+eAOCui0VFUx34ssLoV7dlInIU0GsPedAGqC
b5yGZAuw7298Y9N1czOE40WGoR5pDhwzRJjTpsU7a3zIwqtG8fOj5DkfLvkJfbyR68FbuT78NqOc
6H+EJNeDLKos1FwCzfMcY2slMHCTbu4KFqu6rElnMN8pCtspX9rmxV4zX+SZ/m/QIR901Cx4l2Qw
I8S5bH3qQc5dgX6a0Syf/myCzSsfnH3OmFUGwncsrj6Fw7oFJ9PDZ8de2KuHSNKHrw/Lsve5+ei+
lCMkhUVBszaR/t8y/t2etminyIjgmXnPtKUULFZZAFxpRwj6AZ9FC+E2gx6PkUm74M11xGmpvIq3
DPQsPFlQp6LSM8/gmJxkXJjGHnloKJzpVBltvxnxP54LWq+ZmSxVxD5IheBtVv8aouE9N337X17a
SpAedeGXvtLuVdJM7n09xJVWwdOA9WmcYfj4Nyr+oHaMO2Dg344zNlm4OYVzDYltrO2Wxft0qDsy
44RmRL2sNAgBTutlXPt9VPYqGMFJHsNK3S9TvFwZAeotcd7SnNPO08X9cYoxlq0xGRNHIJbK6kD/
DWQnnOHRJpm0XBVWgedC7mNczbqFhx4gR+SOG16SVJoy6n7ZtBHMExj5BPkUyWEfujY9GV/4Dl5t
YmUw0GP3dfyQQAA2WgQENmsuiwSL5lI5Nuw7SJCnC313jgLa4a3iNvJyFtFnFb7tP8eqwKIpkeTl
aP8Y3U1U2tPxpZItSNgy2z3MZT4FtyWAF1Rvv+1c3jEAxWUwf4qqU9O3+wm3nlYHoqrejJERTHmE
QzpYf5kkmU1dSbRxRTlLyWjcdLvMOsai2D9pQcU4dGAnSv2TKapmsBboXpiAZxejvHdsmD6BaI//
l/xWzAaFX9zn1GKmohsf8zjtBxNa4xXqOP24n4NrS9sBkBSOMHeUZHakXAArjwb/c0+vRlacmNUv
36OtgTdCx/5mEQYJruqvn4k+rOj4v5W5N69QTOSg7aef5nrKgAh8Z5V7Mysd/1YKHcgJfl6mhayR
/cHcdrHgQxC7KBqRjUo0r5LCyh0zV96nCO1+fXU/04qIXPPUzir57Gzynjr1tZfnJWYYr4toic4V
fx2+bdFpTvyUfXIl5n+sLhV83kg9Hxcsy9WlW1FjyfRlyoalAf8TgpUScLsdQRhHxqOIu8lh6YdH
wOUo6Rcz/NTnFFOl48Og64L2L2PkEDlIPz2TQOR2N3L/gJtGMfNibfSDdryr/yJSoLRY1WCmtU4C
ogXZabmQ8Elm3qBnOl+d/RtwwrXf0gHV9vwHgvyNp9qrlDr5Us2598EHEoQTC0awPbBL0SkBdq+T
aT5FfaP4BlNyI5ql8PhmWUJTBZbqckfAgZoayRzWNEahSgay95YQl2+8bMvDdKNZYrLurY1/fGU+
xjkPr9W6s68ymDqPxx4czkxdM+zk4tjc43GKjdtXeefXrnw8NzeWjxxDrziGRt6RraN+jJ5sW4bB
Q33kI9wOXFmdXIx1m3MKY07MY4XGlRpsAUYW0EBXN01OdI+fitpa12ClG2f06n7PcpH5LVdHuzqT
oy07NbY1ThAdXhWAxCeV7dIFxeLUNuPe1tuAlyjV9cBFZ1Oc7s9rzgZEot+wpyOGyP2Y3I1mWcS6
Lj4PYpHPisIMH+kFqUYR61HKQ0lFXyY+s8wPr5JqslYAuBNRx2FTg3BkT2wnN5S7jPKbWTabzknE
A9gOYAsb5JeEM9sDV7LpLJeUfVr2KwQvA74pyHf/sOo6ZDwfZVO5iVEClFiFqOPd2qYbHalW/xP0
lOhaBIuf2aHfyqm2WL9xKaUiDQHRmuUkte6FhqcRCila87U2fuxhIHykflVGmU5SK749khNXkbge
JG5hVNvsG/pg2mlocV9JspC1G2q8Vax1n70dTGVPGJExIkn0nEloRXw4YNHtHoWiqpmoyt4a8eeg
gMAZdPCER3qLk857Y2xwDI1ay2sTKDmtfTmpAeh2MsZiOw2zdgkRNPOARne/MiXlJXJZfwV9Z/K1
gJfW35g4e9q56YHoh+fnIrcqNiTmwG5ZnO8SldMe3XlbuIx8GDqz71xcDH4omBfLcSOeI/FX8N6T
a/kZnKTU2mOjaUERYVUX+dtPIceqX/JYThVIUYrett+vqM+u3kqJmubNQKilfv0Tw6m0Nf4BCOXz
72Si24Zj0HzVN9X8V6S3aV2l94i56tmIrQ/G7T3uXbgW3VRhC19Cej5PeJ5rZYQkT3MwIhiQ/AU8
jHsVE5jtCAWl7gttrOZnCD+sVkB9ah+30fPtcY12N1Zq8Ejkd9lcv9399I+B58XjqT9bkCcQU9CG
x3eBrm9BYSfCX/AvOOVuy0wBZDnuAivOrVo3Vzqq88aASb1TRAJKGnuTb7KC7ZG986bx5KnDxTPr
Ijln43+o633SOWd9Vg5ndteKuwmZGQY58wqGzCmcINmJKRCqMIrqn6O/J6ikXCS1lFRtZmzIIV/f
/kErC0uke0WjfjOB8oBuCCbiUpV4Hr3mPoSaVloEd2sRNa8nls0PSRLF6v88H0IOj3vp4QsYUxfd
XYDnfD/x7/cqXLo8SILuqEBTSoTFg10HtdrcPdSpN2e9GRShMv2pP46zYjusOcA01J/gGV9fdgJw
xfaledz5nA9TjDw997AaSru0hlIxoIdlIZR/ht1UCN/8RS3Vny1B5ZKlxeJnouuSIHgBJ64vxUlw
/FtI3l7hqaoTzdvSfSkwTA1SemGrO2c+XWXLnbz2aoZVUElm36AFGo4nirGaF/3hnxBAf96Ci5kv
bt9AASB33tYg9e7ThrymHJtLt1myw7q2RF43cwgw+XB/q41rqynf/QiwXOJ1jEbtQGGFp1hQdopa
KFbcjDHBN33NGDBYRrwf1gGSdsM7dpgvbfr8unTyv+89trINPOnPlI99lj62HoAVS9FE1H7p4lhj
vNV2oPY8oYgeuAv7N/wWlq/4acoumWtoMVcyRK/rRRh77O7zDbksI94ioeoMbLb4OXHI5Y+CtKyX
ocjtZN/NH7shy0c6eo2RSI910y4PzCfmZFEeonxB5QnkogOLGZR4lqXaxkxlr3A7O76YTAQnbcEX
GRINKWbA9Ub+VpNCEAE5A6qGC1woPur6NZpo9qSbdc836y6f6tiQODe9s4+yxK9nj4XqwoWY3xOD
FKRBH18sQRWGYmuG+atKT0S949AAtXcV8e3jhjorRHpYoUZ/0WtEIYOdH7AqhhpxY+UvbgF5O1CQ
Xfd2nkH3p2b7hE0p6zdk0cr0yF5kDbxFN8vlA+i3zlKoA6GYFgH336pozAMIeYHl5yjZS4JFAp4b
ZfOpGGfkJOru+zlbfY7UyI5Ac6MLe2Xz8lElc0xpCZ0LqJt4jZmtRXUSoQKs0mILaIu6Aq+oUEmn
Rp2R0EiT3fAGWEJodEGC5O7y3ogztPVYGoKtyjun6ZwVDeVcOBPcKRUdNIPYhl1mkUUbkpwnax6D
SrWx335B2eS7I4KuB2KPWB/l0Kq8xkPT8EqEjkB6GM7LOfv/7JJnkLbCg5NRv1Ajn9d3/xNcdXsd
TBO+KCoq9VM5OwRcomVHzsAMbGlnYOsoxgcvex18s9My59lSro50K1vLfqusfxLNqPu2eDkG/9pn
7F3Xy52k0B6whki2LyGoUs50sGZOt0eK5q3XTnAwoyCn+2MGtfViGrX2BAyXlwxQd1tnRURWqGBg
M6dd1aNvn66d4zORmFp8G2fZoLCO4Dpi8lySlgkcvVYTlbWy47XJtICbJNZFZistQCMXweTK1DEI
o8b8n6dSTUV+v+cb3uEUTJEqfDu0i24Ns3Zdf+99vFfuyCpOVHFwxyGR3JCWmSQGaod6/UR19YEu
HjVyb+Y7BNJ+NQjuiNbQLNVsh9hj+BJ+Q93DsP0C6RMphvxUwGNHd+mxqqlTMp+t3ewk0zhhDaC/
NhLYTUdZIQjEJkIIt3D11pd3nncBUHyZQdEXxHUXlFU/EHu6UmUbIJsuvpYRB/EweEMAhZTJBN8U
U1MRNkjSTEtrFUuJyjPJYWgyTVLup5YS/jImTxxE/1pUxnCJCbgukoT6ryeXgJ2/bCdn2bQFwH83
P5vGYU26q3NqxxR3REO1Tgh7vq8MG4I1zlXtyFoFbfvUDIJd+/UR2G0fCskbzo3Cs6L/5+k2ZG9I
YWdnjsWe2E94m6mzce4bEy9fcJ0ophNWcHQ9cUrE+4+MCzY9rkyGtogY3eg2M2NAvgIbeixgVvl5
oBnl3H8WjTvMGBajz3KDbbgYaoU9lS4YRzc9wyrdHU0Pek6lwsFgF+4lQhergHYLr7PhqlRdpCHg
eZWKiZVr0BL9RuM8CIcclNtOXZWwbJH2TTVpsNDyv3gh0uX3v1sWaBagCs1WZzGkvgb4rEOt/Ast
AL0K0OLNplaGjYAtm2Omd0Vp67IDlZQ7K+5RvIu2RhbTIkdqnGNbPti1md2j8TDazEtpk6wXJggZ
FnNGKtwVAFxUo25NjFGsKR4Iwi31Fshq8YO9oXzqkOFJLzHkeQtY0NBvA7nAJSxfRti844AfV/pM
YyLbltgBQLwewXEsYnWIvXQhP5FMb9GMpqSYgQsvX//ckt/AGv4voIt4O5iIjGoMAuPxBjPdZwA1
aOvHj+zxxUf7lQYsSPqQjngSRRkwRc8kNgeW2zlmcUM+jw8iVG74jk3hMeMvId9Lxj2pVXJqx3X1
yjbzwEqR62Cc/OVzvSIk5Z6JAru+V/a94PUReGjLy9fbuB7djICr5I1iWogMbXfgr9ouzqTYEie1
NUYmLYIp1FoRqTp+GV4ZlEup+rM596v0yRLeIN40S7wPU5FVv7UJgXcDwYPIrVb5i4pleD+eEch7
5ZM/3pcajzQiMffWS5ndlPYDDz5xpEBKBYR9ZZXtVcgE5LSJenaf6oRVNYz6OCv96/RmMSguI32I
TPBWBvqNe8uKKcdwsLrNwFz8IvRjmpRkoLSI7aUh6TkKcZ0sq92lbonzPVYHqhZbIhzu8prf0BQ1
sNU/qju9uraRTQ+qwFrxaXiRxzuneNGEsZ9gCHaYtcJM3fKLqx5QlMXu2WvdCdDMFu+V4QnNX8Dw
G9cvQMb0Ncc7RUm084jfkASixDIygh7UUnwTfVXHbdhhunZPqVLgVafRCQlPc2+fL5jJXlAXejiw
iAWr7jQ+SkjwPv2sdBmJGrIXho4y8Hm8jMwgK2mgxwMINhEu99KPrnAbZC8TBIqmZWk3QBRskTIQ
Zm2CdTtGYxS8s5ZOHKNCPnsqYTKS1m70uK2a92yJ8XR2cxbjfCsXRG2EkWVmBKzbi6AJ3rcsOR3k
LjB3lHle8txubH97ICTVDvIvKShoY6JtIwDZQ7o2/MKFZ8DXx8ZaP29hlITP7KjnFChAeDXFU5qY
OCH0ONsCQyg+b87k0ZdPquF8VrclIvPQGXcJV9hnQMf5pDISW5Ywu6cJyUvifZsmdVM4XHoV5xPC
oA/g9gz6dAVxdH2U1qky8/x8S/DNY6OcXAf6wbqM8J+32dzG/85xBQLA3Kvlkmhq8tU6Wz4DTsvQ
mpRrQp8zF4aVfHFfbAVo6j1x6NIpBI1w8PbRrN59MwZi526ZHMcv/EagnW/p1pyIAL4HpOWehT/z
Vkj42y2IzIc3DnMjIvxEqBbe8L9dh5/Q60GQDPSea21gviyyvYstYkmfwcozmbb7K5Nc3fv+buJk
inS8f4ufgbJ7VLDor+clwke4H6QJ/piCrD1e97w7zS5gLxEjQkIo5JiYMqfV6X521dJei2VgCCGE
6vpcd1ceH6HwfyVm9IkFlcS6jh2HQC8w5V4ZZYbFcY5qLevlIJWpXTaV1iL6UdpUm8oFX5v8NnQf
gDEDkMpwUqa8f9MjA0gWIrnvk4A3V/PfmvYl24eD03MN+YT6DF6TzC/CapYntL9Mk9we7/Ho0o1I
IZkiS3knLERCqPl2LAdKqx9oQct3En4zQd2D5wSHsVhvvYbKqwmCTYH0hUW8zjzOpD05C5eLYMX8
hQTXOXQhTMjKyDUluZ5tIyrRFQ0jjDV7QhFuRi9SCIh5/VRWogjf7RHVJRqoqrfaItCZYcphp5aq
BoteWpCh6oD0TvH/RRzePvPeaQugNzOq3AAOG5aHwXByrOuSfJV6NnIlh3SniPnHJzWxPVFFICkF
DQhrKoWrQwxcPlV0A9Cf/Z8+B8HOcsQfZCVio5edA8vxJEuYZrnPaN/uKr2+FT0iLeJlvdZzNMUC
T/mkRxl+vRPsabS5yi1k0VeoqUWy1dCMXHEC1ciVeniBzepEJVkicZec1vqkcPrU8J8v/yXbCkiX
7usBwYty61B7CkbquQaOIF3+vUdo2SuxiRdiOHgr1gcT4xUfS7vxTch0xQEH2zkKl8lNUuSUWeln
/ZPV+Pc5j3nZeeEcHd5Oh1+fWGo56bBr8ZTQy51PbMTmaCEQxwIcPWI4pXNZUlzboySGiBkzyhTi
0Xam/iazMzI4x9qBydRuuWgY307xujaQZywgLXyClKKt7RQUKjJp/Qlg6BIxQ9gIVFqUimV4P0Lm
ufoUM7pUvLjiNEqb9SukAf1TKrNTTpwdRxOPtnylTTH6XdAp3vkp1m+/7uNuU9Lyu+LXiCYBUfda
ysUf5XDspJDlGWveEk4NgKY5bXhojyGmEW1voRogu400DOOnE2iqpUDUi3BFThp87/7Kb+djCkJa
jNu8wRqmAeiK3xS9fwXEXIHw6LWU7yR3oY2GyvC5hxCLg4WC8/PkcWt9ZQFuUFM8s5ZuDn4qyzSF
CEMxNrAa4xpQ0DrgsJVTwzCHWv1QD9KXEgYGE2KLdYP/NPIif6sGBAEr0IMUBOy/Ce8u678FEWAV
RlH1d1TZ9IwvOpGUXGB2iGt48LxVX6SYQdhccvT0SiuJG3lBp2KKeawsTVb4OAwrNzSB0YEZROqC
dpE9Yr00niYsRYmOVeQhyIuCWzeab0ffn6T9JMOmI5LhZV5nlSo9xrEQOHtbnwOODI83AsHK+Jyj
t/iizKJor3JPwgdq1IpUT7ZUgIIf9jvP03dGra8x7rCPhpIdy2cAKk+J/eg/Fg2IbKNGIJXlK5xB
fvnujzrDiYKS26arVroL/lEBFU30EEICSDZk8hVrZ6tfO252GKmZOc3RKt42MjdJJZ3WHVoJoHc4
rZcjr8WOlSoU66g8ZSw4ZdlDpj3i5LGNBhCiA+Y+1oHzLd2tqEVTda1B0wL/QTyczNm2Lebd+mYD
4RWretYyBKcvbuum+M3pTdWMm0lMnas+2CnFgZp7bsrSqXTRpiKZc9i8Jf7h7yuXc9LzjLa0Hzt6
i0W/+zran2OFj9C8tpvN/GuBO0Btv+Sw1YBYGSVw+tBMdrZmiy4OIssskqMMFflH8EO5ypdSK3Wn
86bHsQMjxHMG2jcyFEoC5fZV2p+WFaphJc4EBFxbuT1ZyMcplltnWiDwTjCc2iYLkd+tcgX45dp6
V7LBmdwK7bgcj2RE85ut2c6qh5pM6mEKk39UIaxwSwWiwuIZy5X9/CeU3trakoLxMmy+1Qv/kJut
jQyl2Pn/tyjIyb3FDrRsizKELranehquV8OShYDEjtV9xARNERDr37ExhpXDCZKLw32YD6EfCw+i
QTDhbeQoWvsufVykmew2eoMP8/kyw3I4DMHl+5QdAXmnmFlYfrZzrgAybVFhUKmsLr6SljNMCgnJ
O7BTZ82BQnDMjaNKrcIHWDckOc1cutNJcRWy3FYIRLTZ8BrANkeG1u31h2tVkRUx9gMZjGWwOm6A
83g+VAZlv0C8qbBoVJiYklVDXVAAjM4eBWVChSibeFRh1GgWvVfzA1Y1Y87Ngg6ktEBwwM7/45SE
37NS+MMkWFsdJWBI5rhcW1agPnAy2RbOniM0GjrHBQu5SEYK/YYEO9KUM23e6WBfmez5Okl+EKRb
O+8CYf9qlXHAlU1UUTTn5AfxBJ1Or8n24bn3+zaq55MyjbOyLFCxrUgvA12qcJa4JE24F9V3SjM0
GH0GY6YWhb8+PJ7BZ6VdwilFZmSu7sisoFtUqwWERUy27mObL4pubFlCBEayqNfG5mbvc7W1Xf28
m9Ly2bLx3bwi3vfw9eshpmLeHsXpYdJagFLIG5wlozJ9vuuIYs68bMy4JVjP7HCm00cuskhWWsm6
l/JO5Agy3nMPLahrYifNSxFXzSmVL5rk5pEX6O5pQwQ9wvGDNl+W9mpV7nDYwaPj+H1IjNGjZQhn
8xEze6vGkbLA5l9yijAarUH7843VbXydDLn1iWCnWwzDDM8r0v2YStPxcRt9KFi/6bxqH5LjUpqw
2d7oyccN48A6pQFDkP9s4tune39h5DDzn3QVb5qqRvSxnqDcuSihpex85YXIaYFxjxuG8pVAqtRH
7fSnVmjg0qnKvkdeFaCF2CIWtYnDeRFn6ae3jZq2P5mWxV5r4q+m86f9fq3vKl7EVmHyM81rKCK8
XruG0QJVcJc227ct2RIptCAZCYg8m8rChKIv319b9Y6dEaDlSkAW0bHMQgObdJLjnaepFZHKD6QS
ILtlc/faLhaDjRZ96LvhRlxK2Zc8nRoG6RjsjbgGKiPbD7aPtdTUnbqX/eC/tfLaKqv+h+I62/Ph
5h+ZJ8ciZLPKs+jtv4UYG+UQWtRVHEEeSb5dDAlf8+AUZRK4KlkYT8V7EGd/+8Lyjt0yyPpNkjSq
qJUsKWPDtWdHszi4Wd6KnKeTgOrWlqJGXhHRSgFoNlq8gXLFG8V/yFscuhH6vAXgIpMn/RRLtRmV
I74bW0Q1IFXj1d5gE5KWJRaDfBu985pDjysEoMKL1npZDl7+on31aigEeDC97bfetvB+5lWOduBA
0udoTpN9ImIfgCOYXtoDfcKuoiCQONHKsvX60teE8Clc9yGY/erZZTr3MbYXGFkQqCoVlvAR4Vnz
MarixusIllrMUpMvOPEfD8lPPgQw4sUj9Fjn8S5wT2ccwj9k9i1AgnzIOzRrZoB2nPywPNtVtsrp
fH2UHX848L5ffJdWS+H8AmgX7gtijhsb24e8RPXHwTZlU9Bam3HqXnRXQt5b4cMLHXPZu7wu4yBb
Vp3gy9baqNPQC83v+tXEMRMvYOlQclpWLNn2AMdO69BTuGYC8Sj7Xn9v7ITM23EDEx6MuaIrAOam
AjhGYUEfTc8ftJ4MiP37WMof5IA0vL1Io5HLFEVSQu7dzfh0ieGifLjUrLNt2I/iCI723cWWvQ94
9AuEmaN9+HU9m0GreziHDE/rzodlZl2Ftlx+Brt9QLoN3N7yzqqdppnFmvwrf2oKFb24lop5+9gV
t+FJttT5lYq8qPsf1Xrqdr1MwsuVjZWl5r4Vg4v85QzAoslZkED/Pc9CaLcK91BN5t0lICv5A3Bo
ogXKvBrwZF02WBknVJLzRYcyvkEoTZx8rkMtfHHQtzkgGnFsZ3WwFI/+DXNsZlTWHSPpC9m7Q+5p
OjvHGF8la26RI2zsTmTOyq4tW6qJPbZsLX5DXvd8XaPgRtQOrD4FvYSC7S0GMBslB8fGqUOCPgUf
FZ/OKkBvXpzbErZHgE/9cjrm5/9GcaocBJ0HoEgFopDVOqUXzgP7JFxRA3pVmJcpOydM0AzwSpY9
TswWlaYFB7ic+KDc//tnzEfers3bhGTbJAVPT70ldKAXuDRYDViMDCLGvl0qmRzTAVWpz20hi54w
vvc2S9lvxawcig0uOU6U7isVc4206ZEr6lrZFctwZfUeG8xywz4rri64kfbqOG5b8GdCuWyL9qyT
zJoE6UrIPZwTvokvjeSM11EWn3Axe06l0p3clgyJN0Rw9cngv29RSzR7ujdY0STsGKcQ6ePxd4Uy
HPfMOZ+XBDF6gWh70HKvKzZMhJphzRFuy43Tg4Ejc5rSMJV1sC5YRnYyMCn9V/bWRLiBqC0gZSgn
/KMCQ2mTmWgb0yPo3KjAKH4IERlNbDxTs2teQuO12BUaJ8ZrKO5EYX3muYHFk+VzNVbq7+sCzjf0
eBG/EZb5WDdIzznoD/29zuvit1rawl0idHeRn0nbCSLJ9+nADBN7GZ6milv8K9cFqj4xsOarSKzm
wCVbw8LV/EYBdA7tXFzpIXlap0EuYM43Rbw0VGh+Vph2slj1BjGhpPduSB8DV6a/W1UZNr3IyqeC
gd+zvIOjMW/kGWoaALxfnhMnoviQYxcGqQbnkqjJW3cmL4FbNTCS1xqfOXdvQ1fQ07CU6zrqknrL
C0l71E5UYDOmPM6VCOYnYmkRH0qiK1HXEGV01c2Mve7H0v8awqObV805IK1IERlAS0mN3EH5DsGe
OiD12xITqZIjk5uQr4N9Wv2FBsfZRHi8P2SdcnUMHAzyXP6WInBlXOxywJboM2Kq6oqzmEZSZixI
c2llPiBC0WIQICsNBnahg+8Prl6N6Th2z7argOY1/TKqj33qnqz11kn27uThCkbq4NKBXHKDNSXU
73bEm8IIOhMfrZMVcs5Yu+qhVzuydt+ryVRmTKaWCKKZfIaWRP22WTWQOkbUczmdqEEXsbCzKMJx
vCwcP3QFEMDcqZS4C+dcjsLoqeyLZ6lGJfQa7Ip0YV90eCD1QG20DCasHrrccOq8PfodkAoSdiNz
2Myj8RU8WCKU0UoLrd3h2I08noaakoRAiVZwQfvKQXX61mVfv3Uf/hDnb+C+T6VOaLsyBxNY2yO2
7QBYjU+4vZxmlVIF3cz1QAT73BPk8/a3B30h3a/5pQhqSgGx3OADmPetpJwA1cuYYwTj15WgGOJ9
MWYIKQhs9SKIgYbo/Tlsh1HyPBnHLchrpPB3PDEwJVGbQ9ZFUyRHFj3dKzbzbcz+l9o4KVaTFFr/
qLpY9Y/quGep+DBJJtDO4wcQ7wRpnUjOtkM8RMF80Ctd7S7Kqt4Lz69gUXIck48PEaO1G+jHRaOr
pJmcU6pdJUcDn6thGsNP8knLJvIlnNledfcU6a7gkw0NI2Ykdd6x5u5fDkbtidBDnKKnfIqghfzW
0ghe35DCigbe98d1mXCnVARg/tI0SCN8nPOxr5uyTW2RfqwlSpRNae20KXjykptmtO/0VwUdTYpu
/Msoyqhc1jvIq7Lq8nkK3v8MFjs+Drpv/jYekGdnUfgYqqLQMAa6GKCfj3wHscdMPu7rdg8nI9XX
AmFG9Y5fD6dc9RIUtzVwfopQTZse1YisZtR5fsKjC8NydOl2A9vCmc2vJWLoAWI3rLfn6N4LCpB8
x247U0Hx6ogbut7gndjX1Drh3OscXVnclYNr8KgjqqKaWNTr1DFJ3o0uAXxKmCYWQ2JHy6jeZFV0
5/Ch2T7wTwGYnVvgPTWSODzJwXXETN/J7iXwJ+RDaAxuGtZG5Bivi9GBoZiUKYygkfLEmldGzYI4
+PrBVYA6Zmdm8azZ6jvWO7tPHiP2g0nYCPtiCb4asW1dOWhxkdplJ8g/A/SiX1B9J2wwpWfjjgaj
U4hz7cL/iBPegDt0ehfjbT1bYYhxGpGOXRqIcikJqY0p3F/xw7TpBlpNsR9vj5kD6a/2QsGhcPoh
uLGwR7ReOwlDZO7k00lk80sIOVo9DP/cMFyFd5WBl/jqhRpIB5M1Z7u9QAZsPOVXjpMX7TugaBN9
Au24Ni5I8gS7PqVOkazTTDEMKIQ5QeTYHG9/1DygzNGhH34LRr/gGvsuQTD3kCFGZfxIKKizVDFd
yMTNyqDwoSNjg/78IZ2uW5IaF0TkCQUONkNvvhjkMcHEZWsgdUWny47E8qhJu5NpZI+vfhYPhcvO
OzV/nW1ygOx6HxIcLHSILOAiHPXLS0f462HNgHG6OegEy2qoQb0/a0rKR9cvPJi5WfhIB86PoAf+
Lz1uaQvus7JjlDGYNJf9+K7UEQyzJ00SWNhqrAbfjv22DP6UYf+Z2czY0O/jM6ACICgRGm2hzpTE
BC2hWuJSHt5e6u/ThWEK9yxcV1iFpTTLum2FXN13QUy1INHPfgdI0ma5rV3n5Kf8++sox+DXG4f9
udftL0K+7GMOB15ZKAunXf7Ij+zadVIoBdgZPJ+yHbjC7D52SHVJg61OqK0kXChnroZN/UsJz0o6
pq/QMu8n7KUH8WNczMQ4QNz7tPRyMqu0Ht2vZWOUsch5eq3SKZwn3Oq0XCI56xbrcPwYn0NmkqVR
dcdkmYe57eIZM+4ES3bYNqQGlv13KzyU3cnOvI31aJ64nuHAz0qSMeNdipGJje1Si4+PV3mAelg2
kZ23GaHzgJbVfznTUGilqPEhCMW3ReJkRCKOthJQpf3aE3YwM65X0YlSdZg74LsqeNrTVbSMBlWj
2QtXShjmLVYr7Va9wxZdHM5ToXPVVz5eZ1OyRice1byZKk6WffdLmK/M//M9KfUnpkkfS0r/8Z5N
gmh/5tTEQ20Ui8Qy2UMtgt+/DWP3MFNBVkXEWrBGgMNvV8LPQsk6p8yRVz8/8+qbB02bF8C7vLni
j6umi3X3kVdsx/0PaOyNxLOviFRXbwkUYLE9ogRmt0cJze2Sk21lIpW45Qsu0eeyz27vwyLRRre3
4M4CxDZbiGEZLYx+u4eK8cwwsTovnKTgMG5m5DvYpQvcP4m7A4jJlcOT2Qqvu9O6xLS1Er9gb1lt
8vJQbvxHHasTMi9OP940sQnkp79cuC3tQIpSfQXq3waRZY6QfvDHHNjI99Fc0euXUsDRjUKBVN3F
t07SN2T3ClvMPy5irNwagwyGOdnzbqbG/KdeYTvoyC30Mus/O4WmkrjpyhN2EI3FGfHvz9BlHW/N
+q9tKJ+DIzLyVIFaR2HDN7v8k7Cs6E1NkBjsHeFmVKjInh0IhubSU0JmqNwIqwusvAptCKajr7UG
YtM4SJZ+gr0wJ5X+OM898wlBqP4Dl1OVLkvpLL+Bd28HJkIIVE9QR/CF5Iv/9GuvyXndLfyhLVVH
hI9tnjbT0EqeuO9CU96sJMnC8XKTpIWWtJ0oi7yjUu9AQSQiigmBweullQ1KkJxp+EV2jVljwY6J
cS4SMb2Ira34oeoUtEs/d0qudLjCP23GugahoTgJBNHjDImXJH3hlFuDhTitwmWzHVbI5NO+GQcX
xxj4BDmpixrxSau0Ggk0uJxmYxbCmuiOzL9VVdfhb9QpFGDfvOtZlpKBprDhi2Xjg4hyEMkAPDkp
GLw0+8xzC6HSkMraVfp4Y/MY4zGRRytgtvIYuVpiGawaSj/22GgK0SuVxzy+9aqdtvfnWJvwvnDF
lsWIIMWuM+D7wMQx3LuicD9KmLTgPzqQ6kC5zx+KaP/g+twLa0yAB1gcYsfYsG2khEyiE78/FxgS
U3FHkcraYG550OPUoY0MDCHhDi3ZgGTDUFWjSbGx2b7RjXZMBi5Wuko726EgaoZxwu5P7e3iPl1z
BV0Hvc81Hjp0tzYjBIM85Y3sVn7jrzeNgEyO/L0jtleA7hOZg4yRbYke3ArbShlO6vDfwsUfp3Tr
en4ZsRS60gjHVNn0FItxSCI5ydYmgAUCKIN9kSdwVX40cKCGHIzuKltjK/EQnKyMQUiEWJux3rKm
P4a0ocRN8jJXylR2zx9xY/JBHt7dgK6EpjYPHt4VJPrakqL1/BXehBuV21UvMHt1gIwDNnuPyCQG
N11pPJz9JsUN7zFOsA7IMJI32D8dQDtLyx8ST3wpS+DlKSSutTKZ/oSLBRUnqqvoGSECFAynrhgD
4miaowU0y9FMOR3aAPAkMhYgrZYHWlb6efqs0Y9zJ4wwps4Xcqd71xgJr4Z2WfzClF/7ze1MSlGE
Hw4F98XW89+EbVK+d8yz+epFgijYXwQSuA7pcRckYel2GHJiMQ1FjnOBTmd1T12svAkKem5Uyh01
Lizx6ICJKTTrbskNTnMDYAnpcw4bDf1lTX5JlDuPWO1zfVDCIaeBm9tRIhoCh3jbqf1D/ElJW28R
0vycyHTf8q1f5UPmJPx8Xva6peMQroU/GdpgQzZqTUwt3VMzuFZ4xjXCLbXt4w7pjU244IUF3Xv8
Flw4t2z+PcXFehhE4ATDD7U9sFZwOETeY6wzkHk86iiqYp6Qkd5OtV8QsG5186tob6rTbxXFm24Z
vAgF8MFmJjGDlOtVoJcm9iSZweO0IWXUIA+1emJ4bDb9ezA4TlEf9hlpNggHeQBL4QIqgn/A1g+5
gN3akCjUOZmDeYqWrTwfjeh0yZgqotc+YKijwrJ1MdHnGhM7u/7J504BlCtK+gsc6GT97FT+UMZx
nyI63afSb/CW1JIRNRQSbKXhAiE3z2YmTl740i9LHhFZ+vNsGDHEXm5gHiqSjjk9en5Wv94hPjUa
Tv3aCok0SPUjELsfufTWvdUAHiHW28LIlOj/XBjfiIwQ2P4DFdzTVNAxTMRc1XyZMuOyW9x6WJwZ
DOdc17ovZErvrq2hLHNi4K6/bR8EsFipaugQQKCixoDiVvtmXVyJU+l8trGz+ao0MNqdkpFBYRln
W9rMe7HPgEaNaK+36m0hSqcTlcj1iURTDvIS9AnAYvmqNygle5wgr1hO2/1tEncoKYIvytVy6VB+
7ZVARds0LAkrGAOoemuBoqmHWBI89SVTkDMBYGvXyghoxVXD5De8YcQCUvwe/3tbf2FeTpfS4tdK
qFKqQfTIdnhnpcwma1XfzC0W5cdD1HyBMSUFux1PaNE9nsqwNS73EXEtWT4yC4x1y1oJ0RhNNXZ/
+/McWHr1FABYQDoqdorVXUNdT60Ue5cHH5ueC4Kdr+4PUp1mweN28FD5qmG2ETyJb2FPY1jPEtmT
PzeOJdIYREz6/y3KuOjXQaCpXJTXzA766bAJDrjPq/fYAywBziGsRsBQTKZFLCEE8lB3aoZhyXS6
5nQ7La5f1QSpVla3jzhA9A16gjdtr9gtPFq8jakJk7bXDc9hhTeUl500GAOXLdSQMyvqHQpIObKx
ZCW2VcTaCG+WW3fq7rTdqsw2+puhq823w9o5EY2dyn7yHYPlhzUQXZVJUMc34evJzpONWbWKp1E0
Y2HGG5HeFHyI7Fk2c4qR3SATa1HLn6qkJ/UmGE6dbszhWoujHKRFIuZXtF4Yhtn0CWkX7cASoLyP
f8hGVwW3KDkvA7YH2hjX7yMsOV8fB6vyXF9USiiSaVP99EQRgER6SI1nhI03QACg2KK55HEWo7B7
GLG2zGUm06aONufqPpYFAWs1l7cBOHbv+3iLrsxY0SLFFnHnevLcl73xRmEm/Q7V3rhr8o8M1VyN
oDeyhVpYVBObhFxz+SoApOlXFe0dSECfknUGVUWgC+bfTZGTR3OcDcMEtAYNxWzzNL607FgPiwjt
9gZU+zdQ1FO/O/vgjELUurw0MTYZ1ILh+PHMQ0/ka8/VSfxk+FZTHaMoFcZaS+5AvM85v0bBeHgn
xEi7SBxaTM6CAoeP/BaVGcAdv+xsamiPRYDNOcqsFXgod9fVcDRnxOQnu/es4ENqw9fC7AKdzMQw
2q7GJMU5D6HcEB8L1XJo2O7ME1lUzlZHIaha/TR00mQxk4ytkO+O4M3eQcsa9FUprTfJ6IF1Mxjr
c561oIRIyzKnJw786PhbZc1Y2UOwGzR003UCYPbQSyVXsuELxXyEeSGdz+TvDitxNKzVnRCL3WSj
rU7i3gvNVJOBy8If4p07clNBhK+onH7OrhHDY3rVriizT3F8x7916pNXGj/BzYzYC6CAVnNON8nV
RTa8DXDzjcPeKtkh35EjUtqV5joIKlO8KDPWkkBZZ2jCSKqdClG/ZmUduDhglL1i6FIPxPSA2oOv
hrrbcOXLCOdd2REkEQ6SVunRbmWw4ek3BtuuRL1S270GhcKdc2ySlLcaHdrruNQRbVkP/1UMclOH
ytCdsxsCjNt8mmUT6BNwqasj6MLo8drTDWFJlYIMwK9M5YwA62VaRk7FyUbOpnuPbbaNWN98haTK
CjLUlxIv5z2mHAwlX5ICaWDDXAwygiHXix5XAT3XrW0OLORXFvTIFb2ep3UHe5T2KtVemAYNo+i9
+8IHgBkEcDyVAa/Ps4Ltj1i6jgCI4YDVUkJOAfKlYrRWfuIsyawLahSmqUtwtUQVMPd0hOw+ndbQ
IWJpWf/NU/9m8zWGZfEtiBQUq+O0Y8dv4G4gf0tQff3x03chrq57tfAlv7ros5ZhNbA8EbUPPP/Z
ot/YlGadfDzwvqO6K24QEKjf0fxVG+KRS1Ki8gWXan5GTpDH0w0We7CmrIAdfgReNcydpPd+YAO+
dipyRNC4iq9EVV4a1vvvBbRU2GYh3Uq7YSkbm4esShpovMt1r4LtBx+kX2GJ4BUkPCWU+6tVI75I
JqnpBbObJwJ+5kMxZ+VYwoIzEPNKFhCf8LVUJn5ZVh6nQKTDh+Gswztktrgf7K0CxBQx8ZivJZeG
0oI+YEUe+3duu1sEf/Bf3SGaWadYLX76GSZfNsog99+4MvHRLqoJz+q1oLAf0jbpwDLn3049THXZ
nZo4bb2nRO6G3k/DHpOVwyvfbCXf+pnxyUqrAaStNuyA7nECRH/IsSDztX2eZesPtsromHKI7WeJ
W3eKhMjcHrsnAuJegqEyOMnbexSWIlDwLeJZGE6PPJpv4hZsjTFy8A6xkQXS4UsuSGffGClnauQy
ArpTQUhpjPe92El8+IfUai5GiMziV64i4wiIaSPqd60pGjms7VhfpD6YWYSGx8quVVt3gw7uyxBh
4bxI/4M62QoibN3rnDV+IQQnlp7xyOCAsPtrmrWaQKd5uvo54ncYHNW166aOt30nVQ8M/FkNzlTG
HNsUSt8XUBHIckkp6D3Y/1YAQ1zafJqgFfz5PlNv4ojTLFep45CRdW2mk8Jtym5cfdz8D8/0ABhY
zzw6y7zsMAwRC/q5dMbPYUmmZQ15xPewZE9Rr0BP7FvLZKWoHc1Vq0LEL5kAmocl53tmO0V0rl77
IkR9H/4x8nk3aHnB7BCYNjwClSxi5z4DgtQx1l2YhK6W0GSAhKWhQ38nJn5EVyvmZ94+GyQDGMp2
n6IQD2U5zuQjEWmH47BkijQOMalITfl9Q+fhgalF5GRQgl1nsSVqS6kGjqUbfg2kl2Wj0IKAc/hm
INv9zndOLr5BLUOG6xBtmLZZCC5a5kNvg9aETIX2AZnJuKhppkFGD8P0k6qNHeYCGZP7GjeYMAEN
XiuRjkkD4rBR777+VS+23ov23ORJYovw9Nms9alXaD3HxD3X8MTQHcuPpsq5J8lZLhwKwimuP8ga
K1Wq/+RqS/cSvmC6NVccK9/hoWrE6sOFXn9+uPlnWpTTX2XQrCxgSQECwevB6qqRo/MInEA1qXYq
wmzoCkqeYYsmkyOrC1SK+Y+xs0YBcoUtCVN6SEBGmUvIu3jA68gk98RQO3XIR8KJlMQpEwobVErC
ZJEAOYI6lzK4NiFhCFVPmhnA+v304TiMXhrt/jBKL5sCfzwbcBUePKRahlXV/7+rEoQUmT7teiwD
07sh4pAhh9qxGdMhZT4FjtB8g5p/5iA3cKGrcO/sIo24ZWcmyDWI4OwsYjjizt1g+Q+nCMWaCkJL
YG2V1PRpvDrsg78sk2zzztQ48FXTzpvoBLQE4vy9oomqGzPDnisWB26HhyyfrRQSLRH4l50Tqi3/
Uo3XL5/Yp4Fn1DoQhzzNbcZDGjDFPh5upsRCJn9wcBG7ObdO+MDfJR6h/06YGk4WwFo1hL/msiA7
O+5udZV4LMtJwOkyHGAFR8if1j7zygEYVx2ps6kp3ecibNZAh/oz3a+Iw0yqAV0TCGdig9HtrCOP
AartfFzT7vNwDr6TAoCg7uwwOpnWNp5GXUt8jev9BUebl6VUZYuxbS1XGdSpUw8vhQc12/CtRj9r
7QptPCT6glEIlpY+jFJVUBbZgrLAmoQ6UzGeKlLnqlIDSZx4foiL8yTxin/awG/tKGO90ISZuiRB
dGmKTtmB7oH/z9mKlDrk9zhjto63H19E0QZ4sUzZdroWMyD7ihIT9V7Vo5828I914Bho6DK4dhyG
ugN6BVnIFtB12VP6LZd5YNtN7RZ5iaZBWK1IpYwic97O0Cl/gnGkWC19WKiDlqf0yFCrhYGdFA6E
26NSwo+YcEUtY92QYAEvLFr5d8tLJgYMyVAp+iblS3+bJPAw7fE6NQlFYPDCdMdtMYwIYpF4crK1
GRHGmwZgCvqMO2S01HSdRh50JdvUz75jgOKf0+z9YkbtcLHpwyclPSQJNZKXEdrupeKpR7eoSBUh
DTTFDs39UUp3YLHUVaZoA7pQi/Em6NL2BpV1NF9G5CDpKPczckUqhpZfx73B3L5yDv7uBOQlW7SY
RrBe+DEwQcPvha7mxKGgQkn92/WIX9IbMUiwyg1sBQgyHHl8b8HLHZ3+yS3zJJVhCIIFrLh9ymmc
XAzrbxKbFFoXoD0FAbJzOox6XLCGUa/o0nLKjg+37nbthY62KQI0FQW6/jQGZtLI9Ob61SOLbVho
6Y7/xGTfMWc60q9V2Mn/AEmV4H1O7ZySxcga4a520NbkhMHBa8E1avZoPWKVUE3Qw8swpeUHeCNG
Jl3Qnz1DB4FolSPRhoHegsF+UrApRLRlffDFXbnPNbKi8FxWKChvDh8a0DPST0vItCI3KAzIv3O9
Qjo/yfiZY5AItfZlK5PhYuSZCZZLYxoMfS0I5GwtbkyooAguxljINTrdpg2mVpj/ppfQgdhhTv40
8JILdYT8KOgYq5Vase/yv7czlcnLgjdYEsWry3BR2zlh3SAV9Z47SBzSr23OmjnddqpHzKBEPzM6
H/TPBBoDm1BEN/EWh8Ck5BFjMD8D9cQOXLXrHU4KWda25yqBDYSJ8jR1BDdxEA03XAl2gkQivdiu
mbOxctlLQ6CYJ/eQwxcnJboD7kdGDVb5/5kz+NCnswQCiPfAAUK8aMqpfEulz0hDIeEH7msc0Rnr
CsQfUXGNQ6D44Ny3V/kGcu6Z74c7PQbmsyueHSQ0crOyj2cgCf9hUNBLThFsHmy2T99vdOqRKlWm
lY/Ke8jIrjiGNVmOhbF8Y7vN106zohDWydDlM82BeBYS8URsaN58fDFc6y51AvIlYB72Xu3PbF3w
/RzCntxMV1XGnTXPhI+Y53LRQ8hmEZrH8etc2eMspGSsFrNjPFtn9wzYOAYviH1MT2AayLEhLhq6
KWTMBVPYN4QMiEnGmEUbuJ4PBXLAD7iFucMBTrk2swCatbihxA671FOwcpMHQFuKMnLTYB71WELk
G3ekKyt8fGdmTFcXomW5RS6/nqaJ88l2fbcWa8nu0QAcw9gb/qmTkFybraFsiaroyBTzDb5nuG96
3x17kxKt4NaQPUswygpoGythB+bNe8UAB51K4mjpWNZKp2/PLng0sLcYSiKlE604aVc2jNKTgyaa
qMtKptRwZ3gO/EWFMRMfYu30z5oKbltxmqzj8OytpEUSiFYCPHBouAayVmFvAJh1/7ph55Q/RnPb
VPcDjbv2st1qd8988+sQSWb707Vp0kFnpa8eReJsACXhJoLbBDYoJtOPYGgbOrLrC3rZ2wDF8b00
/dRmqPj+eFExRYl7s29FvkZAPGp8j9clY9lGc7l3OdRDWFG5e+qfGuUidq56OiIs0emmQyqTiDLX
OApGEuOoSIFvvDvAG2Vh7uePLaWUcMSNX/MPtF85/UlzNJeH3GTsFSYNYpK3UIAFUx5BpceXBcg8
1M0VeuK6GueJMAcXGNksWcZfBJeHPUM1+rbaZR1sLutAQ91cSlxnNC8h5kxdA+knHlgut3VPbuEU
eLrfD33rrWjQmXzIJLbvuv2GzYmdhbaTMidbsbHc/oTf9agoxj4enpG043Ha7Vd1qPUkyZbXU/iA
TbaVWZQHB8NCnw1pdgBgB4/+dwPDWqq55enw+IVwh9YLRDPlpAm7n9DesdKF+Q6sHGXw2lLkYOiW
zBnXZ5gXHC9+ze9/jdTHFZl1DTQCzCEiaNfqeVfXxt7u4KHHuFOdJ1PfAr/eAEQBMunOb2rjgkyE
Do0VQ5+5H6EhuuV1Et+VR9/gUg5l3dPKQIBHo4NjMaCEDFRgo99O0FMxGbQsvfepjsi7KW4UWYdf
5jKkdThYq7lzqxocQEnKEPX82WaQHL3Sm1Qou/2jmpSnlfy6IxCRnudQUwWwD21q6fXzuGb3YluK
DRbYAhmrSXHrED6VEgoX91yYISoLhCnwn+3SbV/GpwhupppEzBxCTasqgZdKbx2qA7oFaOYzSDMB
jeUAkA7KAp3W8Zb3w4b3UDjuL3S8KUJQQGJaAWSt1YaOT3knEFxpDQkW1ZRzIg014SvdlZ/sMqcG
LkjOmyd84Gl2c0GRqpYNDAqO66+dPSIY4d7fn8xT9DRS+Ktvf6+unfVxrJXsBYcu6lf2x+X1tRRK
baDEHrAvGVjlW2plpphRcGvmdPpJVIhi5ZRtvp2sWSMKYA9jP6g7JPrYZcV9T9LaYRuL6i1dET5I
PpRD9dxUqgSYBPCcPANnDkhU6w4IzEAmosqdnvKVyAspwZjaBvztT/PADrVKXfT5ceimPrCEojwi
EjaoA8ePxpZRGovXzJonE0tT8i9aHgUjJu0xo4Tkfzzgw3u9nkTI0KNM+IxlxeXPTfqMWk8Q2emV
pAVd+dg7WuV/oB6BIXJ3U8AyiP+AqjiSt4fX98HXJIPE5itcUj3y9EEXRLI7/7Dg9Ytij1Iw7rtd
ONqmZaprbp0usf0sx7CfLN+jtLoL/M+2gXVUBq6keT8VkUehZP0UcOB0ai/hDEsYxiEzj1ut3jAW
J/cMhu0IZVPqwhjtYtBYmS7By+DRYUhdyAdXnls8wO9bHpBdG+mQJLBK25qyBirjEAe50J+rfikN
cHUFcQjz0QiL4aM8wFAczcHM9QHRi3ZQjw3VhWQV2xUb1MEY1Z3bMnBXD1EqVzWiYhr9zRZFEvi2
mAMfMeAOSi7Cp9FrMiqfrL2bs36vuiMdGgBrxoTyKL1Zkh2FrgbUgjLj/1P7H+yNuAGuMsJUrvzW
dqdSySE18m+hi/24pFUlR1E4xgVhMxJ+FpkVBf8y6z2XpMSW2MpW+VryjkCvONsRt48vPPLq2DpF
0/2hefdmTtMYG4pTXGajquNh7VkQglCRoP7Hl81jrUn33K5UDDV4GhHcqvtKpKzbnxfYZQXI2OiI
hHtV5qxoQwVo7CBN6a0QiA09W/JGKvOXhf7QzGlseLlFTVBDj24TLiz7OaF+B0VlXCaKJDiq8YST
I+7D2m4O+V9GHk7QDht0qYichAWefbk8mWDnI+jLRwxlRFmAmIBxhvUONfM/ySh3ouNItHj+fWqU
YZQ2IeBzjZUS+GJpPQa00yznexjnDHAmNP3W4ujbwoSyqQEN7N/P/gYJCfNyCnXz9vC0FB2K2Ye1
4KmiI56UIw+Dix27OWYOBMk5vlso/SDVqiGyv0tir1U2S8g0enG5z0G4cPvbCaoH0nwsBefo6teu
134mCtq3StogFSf3rKeKLg21948WfdrPi8ns7Gek4f1nEI6ZtwDEEyLnOrd01zFD15yevEsksm/z
SBGzHD8ITk2FaROnJIY/vJgox3YZ2Q2FkVYy/7hE0xrVRHL53BEwVBojMtswv/QRSVQvYhzQKuwz
bIMDWzvZKh7nrhrIAJMCpBrEY+bVd1Y+KJ7RyxmeNb89f71N88mJqrWz9JUljY+KO/EmHCGS+gFO
tlKbAPMXRB1huKKGbKyNzWMheN5J4jE7dTRMMIr5QGVUdzloZZ1t84ZH5eJKjOun1M+4YS66W6hJ
eqMAD4+OT5PDzck7YQphbwhVNGIYjLe0wSRojHps2MO7E012fYC/mbLkPQzp6TQ0CnEd+Z0x1U68
aTOUWFeGpmF68ITE6lnXy/kkDtoqhMMCh2djdCtDVHRFxqP9+20KohusraTfGxuxP7JCcJduZ4df
kVf6R+SsjuC/RXEvbe76Ckmgrf62OOGFDcooIjYqnOi89H0Ij8cSqDH7LeI7I1HUn5dChuvZjo2r
VV+UNkVT/yGL180esV1Zfwo0RCXPeRUrtnp9UQR15nkTE2DR6tFhf5vBosCdB3NO04lnuv5RFJs7
zQRIyrT530bVf8aVdZrxQxAIizt6dGcd2LgHOKrbrQLB5C6Qlm9LkjUm/Y+jaPazUJGA7QXaSLN2
XE7goQrpdE4BWttJa+HlAiXotJvCeTxNr8sLLHM+cGnL8PNLPlw1DSpiFOh+CKyDdk3X9db36tm6
AeC8SAzROCzyxobdlTqSYpkKyJTg/awMViuLV/lWAzUuO/OgQpEalOaBmJE7ra6tNzEuRJva1Bv7
WpPn9I945HcKuJyP8jYFaSx1HbVjqWVredH2Uzlhdra09qynI/uv/LL0yeR1OoYQh7noJCsS5rxL
n9Um3HwALxRdtFs5+Gp0/5N8iLF8tJ60YhGLKJyItr08oFScxkzruBdoKUWG81erc+J3eqPPEefa
XDuT/eJmIFkiZKLN+klOQPFldjQMnjIj/OlAmN1CdfRSaES66/XSDbycTIizjr8ZbiG8lKTovUfs
+ngSyogM3HTXALrxNtaNoln617iX0NhGwduJSrH31amVm8t/YR8aCRzT285/UFp0B1zUmLydt+MY
I2Y5CYOYV92jPcVpCcfpG/Sk/ZRUbZn+OSeR0IyZOxhcl+9yNdNOqfC0E/yu9DUpNPmv5uYVT5hz
lmg8joC2BupKBMA9YY0YZ7YIenbVOO9qVTtsjKCLx0i7mKSC32mer31tOzrPgmP4By4YiK+AQrj/
d2o53Vwp8HSrJNsARakO/OaN358gN+H6jpkPGkPEiGdYyDbzBsSVK4XnV4oBjVr6K60QKFxj4t9w
j2CFYQgz5Hx7oRfcCprM5KsWLyvSWrIw0CCJTCMYeF4iDzivArMMTFJoOGAu5QetUjUss72chCGb
Bo5SVorIRSKl87g+pHMc5U4D/Hcpy7TO6zU18JEqOL1Kke13jBROTJRHFEYoWDkN5fJI8ErV9wAI
pUsfPMpQlQMvK/9vXqVS/FJ8PwMruYcq9+Wbh3WHjY0l436XDxvT3F5NzXadG+bjPVxY/XDe6qoN
m7gjTZHxEtBVwMjjQsauh9WBxji7TwhLkk+P5nbcikTYb+MKAXc0vzucaXmjJbhZFSwryUgYK2EB
oa6jQgN+yvgluMvXh4H3MKdjA387OUM5yOVLIX4ICb6oukCsErWVPYlQOI2zxkjkI+elPa/xLD8i
PXY7ZMxZWLA12F/yQobM1QXmjUqlRcQ07RgAl4NVc6Fh8Mu/3M+5Wq8DPolsFmIrcfPAt1oVaEge
1Adsn9W6hGS/UkP0vRPXPI8M4fHS3FjuMRJHT+kDlS64HyXi+kVBQ/eXULEXNiaV8v/nBMhNhuRC
Mp3GVy9oxtbD/WEtiUNrrdzt0tYPYSHApL2FcaXBHEnod6AUP6krceUwzL4bt+lN2ma+mXTL62AI
PXX+SsG7+qAheUCuAB4ReODeN9MsY989+6L8hAjWUPAtxPtvvxwp+QYjipXgEw35+CqTzwZzCkR5
1M8JzFWCf+rywSaMbr35dg02+4dXrAdSjuGJbz6WzR4Ld4t3yAD3LUhj+S8KRR0ftZgmCgQrLT4v
uEVgZAMOT7cRWNupnXJ1nOS+FP1uMOyKpJ9fH/nsr8jktLQ6FDlEQYzMFaU4P0PPcv6FqfoEAK/X
A88hRe6mvXyNwBM2gXLz3YOtw2TvRhqPjI6hm/vZz+UVWlQEyPwTb9X6TEiQJKwnQ3mlkroXnotD
zDaiYCQ3CDj5hQsQbaPkTe2aSy2gDZjWqFu0x97nu6uclpE8oYb7RcG3PNn95wnBEgBfJFPaq7d7
8QBZMYKC6Mpj1clnlJFAJlBiIN7C1rdBZogdDcz2XI4sFkyXMUz5PrL6C1TAHoEI1Am0E2bFALFv
7/1Q4zFToxdgV+JhuxZD0JAOJUr0Zl++BmhyyGXCmnAhkdVL4mRkra8GwK1ODw103D3tDNUUZ5Qr
gRO7kILcTTrm4kZSq9tdY7xxDYlseDBTJK3zaUa/DcagjCZ2IbaHwGYOeQsoNufS+9v7u/+R471S
zpHH1RSvybs8X+bJ5WSB+ZAdSaKI6YUKt5jaqHd+qeby1wntBbB9EN/Cb2eN+KyVogyS/+W7OHfn
A606Jyl7uKYdKQr80/lq38FrUzqzbVBn0cTr+S9rmWsaj8n9OOXVzPNIxjs16GvM4ncp2W4Dam59
704TF6t0580IChmIGkkJh5Ia6qk8Clvun0NmWfkt2XhmYBFJMh/LVFIq3pnWgHTSIp8JBAolUTLR
n6grRBf4uzCA0j2ZH3YGL5loUvXQHhkmVpLpB37/zmUzBL4wRxoKDsPEUeMcjSr3nr6TaN1cddLR
RGdMy9ioUafP+UsBzThpdQGPFHb786X262y5duCSaqfKCFmgz3IQRTv4Rxab63S6PU7307Rxg/2B
Ux6hky8jxfinHNIa3+1ypBGsc3jtU10zq/f/O0ZAbyJ3hsnR4gcmzzSpUDlO5phr0S5FWFTZrt5t
J0tgAkNa0tLk8UniuQihElYDIBOf4ITu736NTL7Dnur+fZBFSVAQQbheQ1EZb7+4PpUQ3TmQXBDV
Sz9d5zdJ3B9wnWz8VyneD1fSgqDE3BsHWPtHH3sF2DA7WKHkLmpKDjR/u73ZaT9ND3FL74qjXW0W
5GNv7/om6nSEjK39YqP5pEyyRL7c6fSRFYTwhVkw/fdNA1GUhMHBlJOYydEJqHz775RCBOa8TjA0
7cTwYRG4fBza5Fnq1DWG0qinuoi14x9uCHPuyVOGqjr004z5TAxm9l6CKr8/bzEl/y3co3CtG3SO
8o9XBFNlQp+lHDNq6ixh/zpXXlqWF8JHM/AIJUjlCzXKVrXifi9zCT2HoL5y6w3UMt5fkITiWgNR
ZmUCz0jtu9sNqAnmFiISCtVycsxk9CJ6ZDdaytgEBFRVRJakeN8z8OZ/07GGw1Q6kNBMbv0tOSTk
4GPs0g4LlbcU3ofnvX7XKWBqdIQx6xpmgOwx00BUON94qRP/uQ9R1KKs64Tq6EaspLRIIHb+1VYr
cI/tljbNFjNqjat0940KvXsqmPpW27rEhrwLMfv0xReq6sLFAd+VKfU34VvBOn4EpASoYpfPCWyk
zQbzUabSa28ujWMcABDHSNPmq7TdmeUyEHFSZvuB/DEXdzSV+WzqqFvKUjrd/d36+lERQ4tXoW8G
4aPsdGUSy48tIZTli8dTMTNXMOYapCfRthmvuGyFFkd5hPgBRWsU0ZsA6JcVVuhg3q99dV7XJbKU
x3ImQrVY37w4uBixu90BlOPW2SfxGoqLAn9npw6w1KlxQ6BAG/wjYJ9/PqYdiTp+xjLzP9Ew4l+Z
aC6iT2P4jDrMZoR65vv/1NuNq9Z2TDCWC2HsyvZXghtSqF6CmNsXKwcl1V95roPZ9c3xPdOW4f5X
v9wRUZQKRhqjy6BQWz4VaCZm9h5OZcFMhnQlHPLR6gsaeO5z9dM4PcmIA7cFQiKvwEE1lbVKLfUq
Y8J/budkGZdcR16o6RdIds6Qj7BQOdZfif1uAJzrdsYlmQfKG9wj6ce4/T4XOi5WtvjRltgN88eW
DClTr53GQijm0fTW97hh7pdtNbyiXP4BYiHNx6TkzMBIHjQ5SqxRTduSKnx4ELCe1y0iCkixrKHI
GHx0xbvJZnBz50ynMFZZSo8QwahO6goInzr7DCoodfGBD9PjZsW7LOjFjLplyT9B3Le2eW2FqYln
jttZrBluNgo3JZUDP3sA0IuepgyscQXI/YNYluCzrvgwx9QEtDVcX4y8yL2cDeJ7ko1tuTV8rM9o
osjvxXpQ+60TfyDcKWC6f/5n/+85bLibyx2U7y7FT1BQoocWdm45XNaxCZu1cXzRIbNzUxhzThYC
R/STW0Mgoh8UFlwHqNKC1DA4NwClOQbrF1cSDlIDGg3gv2xIQY40ANnaP3qW2dZe6biu4RQlWYxb
OQbCo0fzuql59rhITKC8GxlUFb7OyEw9XAUnxv/8MANoxJ2uoiTYZTHeVB1mzMq7yO+4DSA48e7y
64y6NIpVmmj2B4g3NZbXv9ah6SEFHQObx+Qvs3wrPPhgdp3fhE+4hgDJ+yXM1Gt1lzeA3s+cbe3K
I09u9D5lm5SNRj26wQDMoDuRXGCS6HEtspIx//ZQ/2JIForA2rftyFqP/kaSoyeBlavXD0g1kBT6
plXC2uNGBcZXIOCgfkPYFPdxQG/keaxBMAE062WxmYmZqqqP+g1wXFsvL9lluPNatX7nIpBapepa
Wo9lDFfLUsCecySHmOMNkoeN19GOybaR8WONKmVgX5oYdt8yRh5UVfQxyRw18iwxM6mRpJAc1WZv
dmFkFaq2Am55ya9imLcfE5UJuaAC9/lvkTY9PI6wVL+LldbAiYiG5KdPjzZ7Sja4d6dQGp4UmU7m
LS4dyRp5HubbzsCM8GmpGjMxHa4BlREicwBT0hEIQCR/pw0KDq1z1ruwwmtWwDoyUZm3qKLVjie8
M5qdXN/YXJRsstLOQKTwct2VVnKkkT5kd8Gccsu1DdA/9zagH/ztgFfukUKSehhiAyZ7FDtTFMVe
VKiVqTlXTmc0mZXryKa0eECTUAF4Vgk6yDYIqHcLqDttGUitdzp9HBI8Iy98NsuDHPjSVsS4neQF
oP/rFuDW7ZlDS9jcTA3vXfblHxIFBJAjsPNnDFEDpXiTqaesy0KC+DPfAJQOpQVU9xp+dr0lFM5O
fnNT6LjVSneiGOeZ5qlPLw1glW8AZpgt7olnM1WIgFY7D4PFLlAsDKBiq6V/cNPIe+ryWDKUf3IQ
a+cc4s4ou0d1sNP+/wxzFTKOcH5ZjwcyJkLXdHnldvPZYOL4NbiXIGY9YwFWVLEDKsfH1kD2TO9H
/J3hXvJLdOrV6kVgh+rM61wf7cfDoAL0UlE2nhflRGSwBl5eAarApfhECua6zSIi4egsGwQODrhx
O4PzSNGOg3GQFo9htsoIlA98wRcVB1EjqtQh45z3dAVLMiLF0mb4qcGDJKS/lTiU3n1+OGtGfNT4
KUZurLwXVk4fqFIegmjtE0eGVvstqOJMcb2OrE+EJ1L1TTfjIoPW93hXuSz5cT/bt4t5Cv6+R+Sc
F1r9i9WLmgb/bQn7BDX9HUsk9TThZYc/r7kz/MmSG+AWJqoljPHnfsNuSEaQElO+eNiSKCoFJoFX
q+xk9UM4ryTX2M+nFDXtv6qaGsoYTyoFKkPYLiMvs6eDvOfNchTpHzXfzZDjYLC3+63FVBRMTx6C
ZQzoVHuwA7rq/UbF+cAcHzSFGK1iNYRzWpkJG0HQdDWM0Vj2AyPoYkbWDUaYUUxVS6+csCEHvj25
sxGC/45bTM50T9bMx5zy9ZVfhfs3OwdtjkyYoUK7ey76te2gQnniSaDUZufE4ZpJ6GUs9S0BZevV
OqX9bEvoshl15iudxseO/HKHEjzuuIsC6SclyeUBaQajIf6FD7fsse3yyd6wYgTvHkd+50bWJXEU
vzQVwE1/GgoGyPk9q3SVuTmCYTtkHybNtHMpFsOmS3Wto0R/fRf4Bj+zqD0C7W+V+xu1tmOChAMv
y58dBiT8qlXZLNLODNDBQx+EYMSw88m9tonMYuxT2v2yTizUWTwXMb9zUNhAmZlpS5lPhwItw6Ut
WaScPqkPd6PcBXYwwbNdcVlIk96pS//KmE7xGNZnkCoNIKnsLMnzVRoahblr9Ho6DwDWlY5gAlK9
x61+byfgdOZq9KjeAP8AD2Ri+TakJhvuVXh8Fb4RqLQs/CEA8ljciMHoOUJJawu7RnlNhn2IyKyn
e4etFzJXrLn8ETma4+B7y6jsPZ09CiGFWjnS4xNVbUk50dpvIvgP0b5a8LKAEuHfgY957tnYTls8
7SUqF9r9zbd/a8Hdp0KBi2fOUH++j2ldm1kz9lixVmKRp1MVEc2B8v7uFe2pDHkSNX3LH9gB8N1T
YHcvt1c29NwrFiOgmWjTon8ri1pMignaQCTE+Y6r50COxii46IjoEbeigSQAe19LG2DWAVPQg4yj
AoYVxU8khL7nQ0JKUpvXS00TI0Lz3sOfalHcFnp+NThXIBsywos+DI3AWDcmwZX4tIKAHXZtu4wM
jg0smTMOE3797v3BidmFt8Usq7oExbsfptxogHNqxBikSXo4NQMBFLQeoHqLtKmNZCcUZ41GHO6a
7bqwn2xmZdUxFQ/tPeOSih606qp7cRGb9z7h113NRckxacLXCjtZwj4KulMBnlWbQ2L8D/Ibt1Oe
2kKTN8+U23jaMI2J5zpHJoWNXHzydmPI1rYN99f9lkNNgePtNyUAtvypoLyBsaRft1LddYWIyU41
8vUgQznGH3AR1jR99DhiUbVG7geNO0HlxBOwpfpYcKCu57G4sOVh6GXjoF5nsv6BJz/PfxUT9vMR
1zdLQJTn7XQhXmiNh+udtC6AWz29p8TPTw4X8KZ9jqUUE5svSB47csk289ACirLcfv2UGx7XTbBj
XEhvQRv2keModK2BC5yMMqBv46VWYUaHKmJXroNtf41D7elk+DLrmRqFh8J9cLtnqV+LKzzvFXL+
oR60QTLUdra+uLsgG+KAQtCFdzVIthaP7/XoNOfhfoohn1qUgLYSmhva/C1Xl/n6dzdY9JxUeBHC
ABs/ylHCneyg02R6dmLANvKi5h+uIWNzKlkFJ4v722PJ23/prcH5iZjEQhQi8kFsLSt9UMokhTXJ
/imrtYwBpIBwVHigdi3APbu/wjIOeDATtC+4ocI/XGX5zf/HQeVC2MYG1cnNZDV/loUvWxrA2TsN
JiUzeRz6868wmuLgeHqa/o981LuZkEsZdjVyFpiBJJQUKuCQaRGr2ThPVYYedIUkkX+RN+5diDuK
8nz/+672bMKaF49BjaT0n4uqiqah2Qj1RcpZaM1a0wdFa54y99NfQgd1AxE4VmYsd4KGN2D7wf74
SpCo4rZ1CtcD9YMYmkOYcpHT8M0XJ9UBMOSOt/EbOQAnEF4TQfmYG3STUCYSWxVrJVbt5n4xp9Ba
X0wk5svegO+ctJMncPS6EaEeii3hk4GiA/xCJDN+Gs5hOYrxAbI4lmsvyMJk/n+ippde3QFwDqlc
vrT7zp5A4t74hD+FLZ3yznT0XwhSv1XwST6vRIl+eVtOiGEV97BG+opAx/6KVZlB37WKZjx+v/TH
1xFtEB+xzLepI+pmTKMmsjCsTMh2QTdh8hSAjnLijT6gn9mRel6+D1ofefMdYl+KvLoDBVltOjRV
ejrXNOsfFu6/LIcvkCS4qmc5ujefOR+vOW0uvP3FzPeEz2BIEns0F5+TiN5bBdWChIljrdBR6rOf
4XH+Yx2mG6ffy1j2ldBdpjNjw6r11g9/MgZHKmZIcfcxIRLskL6EU37tLUlCiKdNTuulXw2pPQId
KSrjOjfcUUX3zUVxIDMkQv+ZBXGXdriWgMzxm78rqFEC4waDLm2LmGbntXJ61mRdmC3TsPluPrKP
Xwdm67dOwp65tQX97fChajP2Gb0TlcZtgah0oK2Mu/64ShFmFdsqz9GUG98r6ucydOv8uonvSKG2
D94nHClSKJIdmqyE2FnAhye1d8JdPG/qaHiEt1RoZ0OiSxQ4XzS9jkJf+BnKsy3AAYbv+ycayfib
B0q2WpXo165ncVXMcZ0JgCPDLc1vPqwfDye3v6854ZYawGpnvTB+5uF3N0ivxYJVoa5bmfRb/flA
SHVDm8YQqd0eV1VaopNYbJGalXfyB/K9fC+KvVhZttHARH0DMLWSlu2PFOLvQPL552kHI705/diO
46zIwalGtM65SeIoSH5AycP3HZD7uPz71WpE6OcLHvdIpEBV7m/FTeRQcByKaoCESSSIcWrCTyrD
lOvxS9xaEdD8n40/apiWsUoxKq3073PPUmngS4S+9Hwb0tJG64vHCJz31QSVdb8Tu/3iRrU2VNMK
8p/KYsEYQJr9QgRtJHiWrPc8i0/BreLgDe6Kowd7MVABrdxN0U6zQHQEcOKQFldIhQ8MCRNA1ykP
9T5P7LAtgdT6T0DrsNPjinFBXuMh23/uOfHpTvs+NmB8JGr1eUCkZEkIjQ7Dq4l8HR3A/a6Z5Ex4
EPQ2mkQ5fs6LCfFmuLbQ2qxwpfrJK5NNcFzXvlcK6oy0YZPLHfSDRtpVdas5myE+bLpCYHBYHXY8
41Ov2z0JTQAqoEOntsFLMVkU9chmHvcxMHyQKIkodFA7ktx7YxuRc9ZFnFy+pmdciblALLa8b/HO
GJS4DHE8zABZL4/KFKaNCaELJdp57jaO4wBwP8ath3gyZuIK5RzoHZDlqc7LodQ/JXDtCqxqdZEJ
qn4I4DF8CRzQqYi38ocI8wKLYouFrseR0VLItbNWcmEsOwq2u9zTW77+o7nN3gH3j85UNMNIOr5+
1s6gBBumJgBMZ3tkm85MOURXXprBiUO/DhIyGD9uj/RL++fzLQIJfpX6q+0kwwdpG/dp5FmtXwsv
n0WBh+KgesVP9O7k5FsGEqQ4ECojOpBgyxmCBfYGRGenN1v4S6y3PIP6C36XPlGbT0EouG1Hh6kl
ANuamB4kmxcUeUrFguImKIVPQolUBoqwMSDnGhNkYQWVkTzyDc/jo9RR7b8b4nZRYy6wDxIRpwhW
bg3eVwyhTxExKKEiOU/pLbRjoSr/ibA2M7lPX4zIRvTIoHybNdKwssJ9/7zC5aF23voa9za2e1tU
lIMqvwZOEP+412mqmq2q1MMP2FzUtM4UZcz8F+07BjnL7s1AAMNNaZoHQF4YYDVIoTpmYOuT3srx
ugwLZBefmFEw1N3Hcj8ghAd0H3GWqgdMkiFCxIstO/eLVqjX/wiZqPf43S63ZqO2s0OM1J+MwSIl
Kk8NqOWtIkqZe7M9R/dhJxyRGyHRZ/GhzTbxJZ4aamsI/nhHjBfxOikICopjgU8ypNkzlbMNjWQM
T0CCbpBNP01HH/8G6ixfy5ZxnwHZc0x3gQhwawxEVu66v1ZCDB8b3hWFcSuklQpr78vHkhBKPXbN
tvv8GvAIL/BWE4wCQLjCqJV2vxNEGy9xlVMt2D0h0ic2aIkQ3bSyygWhiLmLaPJ/9IkrGzzxQvpf
cwiG5WfRwajdPfnVUf++LuxZFQTr/l81C31ALTW/c0/xkDwTeasGJ5xCpYyDiGu4y85B2240Lh2W
Fj7ZFPkNwVDDClV3PdpDNVwhnqrj4HzvRsL7tCAuKyIX9OPJWV3Fg6q7GVIp2xyRIyLEQok4AvEs
0AHeaP1NwLNBdhNDZASGKtIi7MLGoQPzXE0/+Jk46G7wqvq2SUFWZyKIwUEyX/CtswlpfHZukn/X
IRYEM0NJKmU/jvLpsy5wRUyPgt+mCzee6fdO4z0QImHS/AT/gwrJW+EzN7BHnvgVw4NhsZGh69/v
nIGZehajUoA4emE+gjkqn3CXDA3qF7B3AbHPh6aaq577OyB1dqISr+dkZ2nzwl1DRHGL0ThefiaJ
7Gut722XD/lX4LKF4RZpJxcSZnvc2XOxi7vhlO/TSuiaOYfbQM0nvhU1vpalhHMKGiGDzyZCUlco
FpS6kJnOr3KO7GN2plIR1ylbMOIxSctNiggN54Cc4vz5f7kQHYu5q9sA3As6a2oGM6vFAGMPAFCf
eZNWbnJAqhMxK1UqbGjZcBhKtrOYPpJ+tigIJmKzvaDlCO8Y31O75luQCybSqFW7x/iMtfj33On/
929Ao+80tOAmvDiI4iwHnQdS3G1iA7GjvnJNr+h7mkpCzVQmpgVkOJruCzCa/a7hx3szpEyS0nKg
htaW569jVAJApgmuB7IumPTkfXTyHFRyrsKXCUuyDayzhzljtjm9oQGH9C/HZoIbHjzyqEh1bBV+
yJV1i5eGp/kL4wSPQGQaMvcGSaUz6OPsq7DT1usx1Xvsn21MBthqKar4Uh/TNq4f91WQ8os+x/UX
a360uOorjuQjEXLtFwZaKFTTuy4M3XFCoL9W7pUjP4s2w9QsR+KN/bK4ZMRADZxtjU8cJPySnN0Q
hHYY0iR6/x3JW7fVpubVtVyFLrJ4blKDEkcT40eB9ts6EsiI9R+qtrw8ZcqaZrdhw5yqxSnDZXVc
5o1DxBLvqmKUYg8HypNk1pSm/upI4YggvlLQzeCssCVgQGuXXjlj6OBVgMg5ELhp+U/ddztrTiCv
zd7n2KExcSfKGoBDfrLc+N6XB1ta8FDfJDAO8O5pCZYCuJyxBWm+r4qARjPI3UoPBEMTBHaSCzJE
KW7dOU1TMWiwx/ogli6TbSsvUZKYhkqtEP5mcuv1kEjp+STzNs18n9v+/1HUuhLKJQOy+2EL6TvF
d7Ds7xvTO3kPG87TBojEtdg08TSPIv1gUVZd4KlraKYoqLqwan/ZEfW2ItaIy66tz4SziQHveD8U
iG9grVXg2I4eel3dilL8deK5rLWnSjLRQc9g+OGVS9o3kpS9ZF9EUUyu2pAGmKcu1yiNvGK1i6Rf
YWTmQJTDg+4QWUKgFkWY3gRcQIMFeV6V3Po57pBLuzYnMK8vrmUkRWsQHrJe44cVx6gaP/esFgev
Lv6LZ+nv4H7RAgLMg2xPk3/iUjeSY9wbDwwD5qRg9EsGZTEJdACa5bcTpITnuYHIoDjzYmAeFOKJ
ySVGmGU8YnYaWnNr7vRUU5H47xmaIGIarfAMID23PeFhGxhsrOqnVdpiTY7eHmwk80HEiR+OFe5Q
JUJhpG6kN8jd+uy/M6bRmZIigUmiURCfmQctWTVBtl3LbonbPXqN2gx1QXk3r4XS6MswYONTm+Sr
unJwDmhF2xV7GROj9HeVBRpZkkZRiEfyPmBS2pTWgNPYEAT4tU1d0F++05cabKWyn71741mZsBHO
YgZ8ZqV8ffVVGgmX+11jxGHSy3C9NdMppuQFNvVbC2NZEGVVYYy2lesD1BELXu9XWiEQhdqYk8AP
lMva5QAltFKG+LWvS6WcMsGGhhC4HaGz4+Kemt6+GjbfPxayPgZOXyUrKDSLhzZOLJ0TkrGRNclh
52HKv5Oug3O4DBHMxM9Eb0AI0/czMKh7WmDGp/QSX5Q0bt03I79WUrktTdras4LFOCdtTsub5klV
gIc0+RXcT5LUnnhrPrj9AVtROQL64pRWGQoIcM3BsyT1xxBxPHf1XYkCIdjlF6+u3Fin73MzYVe6
KRTugfvNHmHCC9SZ1nVKr8i1fhWAGDBbOv9F+mngndMOxHZ2tZGEym1KhK590esqzPGCd/ECdMAe
BxC90GASBNSjPlc3nEQgidBqQY/B6KBGKNRpqp0lF/ZaBZglqPWt+avhQixlxvqCh7Oo2rC4TVi0
gVXAm/9WXqmqxOwt/AFNMRDuzbsNNUN0RgKl+LQUJRP9VBANAbu+Mg/6ITxnGKUb+f+c6/QBeUG1
9EP3F7KM5MXlhpskMvbLrtF12OW4JxBsfLvbZNOLOxtm9SF3OqoMabp6Ic5Z4V4HUiJDbooblGcl
qmv1y8gxQkCAJyoGWC1VoCxYyE86MDFxTQGXzD/jwzVBS+jXgMBs2Eo9EtC0dCPXuQXlMPCNM3xf
H0H9AdcYINkLmo/I/wo3VVSofM10S3/vR/3AF4i/fIo24/B16U1QhoMJ4o721qSeISK0MJTX6j+0
pwkpR+h+yKvUysosJy60gNVQ+PK7QIIdF3v29VR7eYSv5a7grwSZRwapfc2KSzlxZbuwo5IBgS4+
RNFcIt4c5vGmnJRSy+lzoN59skZO9EXZJk2vONnTN8j3FFlGqD9Fcm8Y04sqWgjW+rMIr+Ny8Uj+
vFGtOq86rtECqA0jFxz/o+dsOeU+znmbSEc6guPscF94A7rArKSla8aK2vqBVtNAfAq+JxQMYAY6
xdwNuJbWHjwSwFVE1UKhB6MpjKnO7Tf2G8QwRznm1MKh3oT62TzqHxxHWBamBB/4xYbsDq4ohnSL
MVZyyVJHc6p+lVVq5dYJO0j37hXnJyp1EIOFw86ePbZaEfLK9U69/VRgwBeuaeNVXtQpCiXwfEPH
aAUh3LRVevgsbDNJDIlRefgJfhjw/y96+z4SL0luiKT9rCHKb+/b++aqOTPGEebIypsOuRT10qn2
/iHcBB2TKNFFzNd78Syf6VGpmQ/hZqwtJ+bNE+Way4gEcKopRr2fcBnJGjWbIpoPvtVmITvrOY5f
zQEmAhNm7NOACeuX4++LqU36etz+m4X9xrHsLtUpR45KYsOAZQt7T+oJNx8S7iBFYAWD2geo73bu
KviVfBZerWabRitlb+5zNreoIY7Ojny/pdhJt9qfYiU/2vV2NFfSnWGGQ9/vSiKoSWM/e89s/f/+
8LHLUCtskO88rJMmR2d3Zgq9Gf6ylheQ68mBg291Z3H6sMdqazjp274zi6oyfq6dH7Kb5b1GMcyu
H9YevitL4bcsb8+TLqMyOD0jycxhn5FMry5qlJcj2Rii6BG42Zs86xBRbppWGxK6o56mNTByrTOs
qEiAsPaxqXRJODCD5mbkb0HKi8Xka16gvU/BAkuGixyDUNU3SsFmWSZljmJ08daoAuiVRuOivLhW
tINWf+qIfzAn4rNtn1WVc+WS3+fy1btZ5DM0rHRkrUJLbMtY3ec8H2ANvI7805JWwUz9sNd+FJDW
Ht2RGI40TaymL4/1EIA3oX6OgIPOrn4G8cd1/yvGOTOPq7KvQGWCP5KxCjAlyWa1dgCLiY64fUJK
3bUDrEqzXOB5ZQCLLUUrO/aaV8opDlBcRyeXi1EOiSoLTtW6JbQ9PbfWqt3L2mTr8KdtinbynUhu
i2bt00lgGbCaIlrYs7ZtLDniVLHCTyVJvEzhdqQwEX4QjIrwBts52cFUS7NHIRfL+h7m3gJUzTtY
gIqpJLI0LPc7PilZtIFkqPp/7/2QI/yubCNONFMlQZp3PIXFCyzLc/jeP1tV/H9sGqyORQEBaCK8
eoQ9gaIDZ36TtG4d4l5bEiOHiwcu+7sL3rIcs1pczM18FKOAw2EDT+mxF51qKNr0eTVGyuxJaU3C
C6LQ8iG524XCrCZui4WeXYN9Gk5K1HrdBJufsuETIAVFLKZ2SEi+rjdFilQFibvcx16Qg5mAXedE
LlHw2vO6UG7ICBr0unqYdQ/EuRxTnTb+sm4M1+Ws9OeuW8nJ9wNoLStREPqVIQZUV7heFuElaobn
+53NCiVAPocMGhNGu1wQQcdVVWM0r3t8F2WONlB+fIqL2HEMUx/pccAp5IgqvLEry8JLOUtSWa3L
95h1tt4AZqTTr8S4lLZjz9n+WZH6fyYtu7v/V3ABOgdchHfU5g6d9lozEd4i3lu5xoiBtQcMneSB
KYtsS3jk6EQbpQc5bm9WDGaFI+rjAZ+ZC8OrxbgopTMMMx4eoyrmeFN8A7J0TuLgH0ChJ/eZXtl8
wDlzKQJIoqx6883WG4WwmgsYHq8VvY481keCipKGdSaD6yGDBHdIpFYOx5H1aQ3OrjmLy67sOzba
F2SuKYfjti5e1DeVp5WA7Fh3VMjU8iS/RQTvTzI76Jaeth8XbvNP2FQTNnGqho7fLE3Mokttt7ik
Cr9DoCV3+pDlYX3UY7wGK641WI8xVXiC7aNmMXr3DbwX9rk8omm743upwQE1lmOf9cLuV/parUGL
WdlGgClAUtjKd5xxRn87cpiXvOSkOWdcD4BUD9fXNsZT+hi0f8N5AvtDcFmEYCDjwpq9WqdCBjgs
QszGV46V7XwZFxmpWWU+uqGIlBGAxqt9HUCJVzuhVbxQrpyNstEKCAb5aDpGLj6oHeUWqcQQLh12
rVRpg1R4nGreMcEr3AUzEcBfvKuf0RdCkwKO6Kz9ycVhi9gVHw0k09kLaPfIuW4jNGzSuwO5m0Eg
owxM6EtTUtud7YOtNXZRPzOAmRX2peynIY7PvRnCmMqKg1cJm4yLjMBGYAxPqtW/6vASWIjXXdia
Z75ckhu8lvwy/ZyGxopVcIe8YAAiNJ6Mzf0Qou0iSqngKH4MLB4fChgPCe9/ZcwjnW/eR8aCqWNB
BGzyRqZKrMsK3y0Wl2zPDaa5p7vFW1ByOSS+fJH3GK9/CKmkwrpcNy4S52o4Cpk4j2OLUXkRfKsP
kvOy2Bf5xM+2UbUhUauMhmL5AzGfCFkzENtMapanNqe2b+zY3hvcbNdDGNfxC+2MqG90BbZPNFB0
vveFRYTOh6h6odrG2Ixj/Kj89YCMkDrEgwPHHtG3MiT70fvdkkLjnLg4XWwpIA+b+UQwNciUjDs/
mb6sppHqDwRaJtxLnF/tIuZqp4UcHUBbREmThAR9tEKoKV47iiYZTb9458N7MZYjCoUri3RdYnvp
Vuf20aMk09nHkwPOItYt8Si4sryKpwrA9+AgCTCKkwDrWdfFmyp0I40FwC0s8DzlFaIpqqzSxiDK
L5qIDYIhW/KnegBjJtXO6eoAwoGjIsGONSZmYT/saX/JHDeJDuWNTXxGamED4lhQodGGytC2K2JI
Jll/H/FQHmt+bxy7EbaRN4fTx492YwPmgMQrqqGCnRJvAQ46pfT45JpI1puE5BRblqgf1Md3nUi+
rYOxS/dHGN5uKZ8IPRXzKhm11leNxYgUwYZlPLEemtzOkDRwC8uCN1SyQ7JHO0JAzmAIhihQLoSA
FmstcF+ordyFNB/dkP/GBOu05lBhEAGxaPaW/xBM3OD7dwwiYHxSNFNKE9IoqM6IzjJ3d/dhcVv5
3zfQRUHyfb5RLrOEfJSG6HX4diZfdWee2Y/DPxFyo3VTlF9znYoTTHqQJrbwoZZsgFyAlPT1ccMq
6k0D+eWB0IGttO+XMO4ek8CsoORgerz9o/m5pMCgece7Pg/0PxuxunvzYHqp5pX2xWhrApKA+d8/
LzvvlQOQG9WUjZBPdgLWGKZ0iFv9y+n39TjPV6Y9mt0enBEUr1GFL09ycNW3u26S5YyRilJygdNI
hrPh+f8cexvKyz6AbsJO/whQmrcwKtwsUZj94tNcDyGYySTLC9f0Te0S1GrsU7z+clJ0GlnSpRQX
htPk2BCmv5hC7GN5zILD2gPo+AiDFpAyGormmLfrEVhTj0LzCdbJ4ZXrjGx5r2m9uNce0dissj8g
wQxrgvKU2V+v9TcVNXmldYmbPMAtWaGOOpbu+jlBRn4b3IdmUEbW0oQmA6S938eYTrtSWDSm0JHx
MIgSV8D3VOjX6Tb0TlN+lJVIEMuwI5VDJrIDKLABNCn0UN5MGOPVEhl+kIwG6Pg4cMaBECTionBL
sUtasICXQEW3a04ScSZ0mGpnsDS4qtszEusVsBJAbCKH3Uy0epJQy//Wgv7ERifsqMVSYNQTBIVA
A/Fg9MrTb91t8EaRn3Z3798B+ov2HFAT7t5+Nqoer6MOk34a0Im2q9d92MKWiFT5KNHL8JkW0JBv
NY/NxpSrb3WyPDQ2vOTi8EqqzpHjFYsJj2QJc3pTSCbqsVmGlHH/VkExDTBrjh072/f76DezHFGP
MiU3isz3mOXo5VsHV/cxoeOoyY7ePBCL5ikOVcwPru5iNxmRpm0je7RrTWLNzjtNm5s5cFFosnO3
uYMDAVLJ+Iv13x6NwgXoC1rOgWOCfKbZ/87i8IpYwqeD8MYTlpTAq8MvxZdgkIN4J5i0IryT1E3I
Scy3V/3TNbVqYiObbcIfUh1sHpRO+ZDuOYdUDkOtJqu1nYVAAHNG5sPwv1n7vJbY963uQCxOSrSo
eJT3jr6PNdNLibLCqd8mqhO/YsrchrnSomqIGbY0HrdQ80WIlWQQrOmqY21NS3pme/EBOAEatB39
4kMryUxjgMdts956EfTo6ARiiI0H7vv8WhqojQDiWEuQnY5yY4r6+6T6dg13zVLJRXBKaWuJF5PR
MZtTuYZN+WBfIYRWoow6MOdQ3noDHhGKOgKc4LWJnD00YscpzC54AOsoTE7cL29PcTfbIBi/KPsf
ft5tkWl57IUmZf8WeAfKAOE/3BCLJkhDImcErvvCYncIYHiAzmZhnU2YYhi+kj4VGIjG0/JdddF+
bGtmqnLLUZLGvxipMj3jXgLneql7ZgOBa9G4nBKgN9IhtDvGbd3xXodKOhJ4NChhe5nUd81894hm
UYh0mMaIT+QMLXenWLDFcKiB1GBxpyA2G/WGp3AUYc9kmY8ngRVitQ/8mz1rNF+sbm2O8bOxnEdB
a5NhK5k68QgNnHyeHGKMIWWhOv48P9Tz0y6jKkNg84wBg8ksh/xowOYIMC1CqWj1nJa3A5K2tQU3
G9+bIVoJr02SKAk9D996szl4soAGexnDi4pN81DKa6X5DhtTE6ZP0ugIMKOfFCJe7+/25XXm9LR6
LhWsmjD3d9dsWHVIoVwLTNqxwFiXDKOGNMEBRtDred8yTayoBjnvcL+ymqwW0LuDnkb/qM0DbfEq
yb/c4xzwMC8iyyrNGZWL/1baqTkz1V6bmJ5/BWvy7Eaiziq090BT/fm2+WdwY0Jd+AGDGB2mKC8W
8/v+GEjegGXlE6CRTj3NK17LIcZXgnYEYsHHV1JyVGasvo1m463e4GoPTYaRUtUgbeLTjau9s7PA
f04YFGyNiIjMYb2dkbJfdKrhec/O3Y4UzzcxAzhweDj5wgjsnQq1MxSQxzM/i4yXcOvMUtcOFu2L
OP/F/Bv8r/jzCE8Xv6l7vrxTpA03AjM+sU5xDVUsPx2hAp68a78HKgie016jian2ynxoG4RqENxX
avoGOB8DLt7Kqy6QY6YjA5dOLDb8U5u6FMXa1wOpWdmEd1PW6wSKfWZhmE88W7gTO/9xDijg5Loa
19Beopy/XBUW6f+D32cU9G/RufOKt3zealKaeoRkoK8UD8dvmXzS4B9j08Up+9guNjiQk0SiwMFz
5YXmZSkAm/zEdGhKK/bnHiEUhvFwAFvXa8/+z7HArvA6SK6JkbU8/ZG2D1WtAdicT4mccJ9aZkaZ
iifwXw3TfJhk3couyjEQHeIfSBToEDZUHyv1Jyu/eHTPPJSGbQ4/o8J31IFbCuJ7Ej7RLx7d+i7b
KEGOpBB9D5iy/rzGG7BpmLhViAW3mzbaevh3kV/RZlxQMQlSJM6fkAUHnwhfQ9Kyd7NHyyT0x6iY
2jX8DMDs4uSViZnWyZ2pIspCqAhTyXu6b4tilfeI8gw3Yub9L5b2rZjdP5h28NbMkEPR2213AfST
grZa24SSpDVdL3ZscjdwX0NxEpf/Vop3MlScHAGX9Gyx6xtk+dAB+MxYSDXZSIX6fZu/AVWNYuSJ
kSZXlYX5PwQIHB5P7XrHmyqW4DdJ4GoQRx2ezIapjeX7LxqfP0MPaq0iyyTL2wJuFRPNFZb91Od9
cN44PGF48zi0fNLdTkdfBRI/OxeJEzkiLR09GzkdrsfKldHxXWVyg/Lm7pLEqz5HmWbvoV1aFQ8v
STkCp54CwMt95oWiztB5+tSLlgL3ooJ/i1Prp5gkykxGTc1AD9gQ96uh/k4y51pTtDoZYtfQ+Wqh
nArOJ8krpI9+UBuAfGKS+C5hia40IpeOlfNQ2YoIQn6N1utCw1p1X4hqWZ+u8/XLgX7U4RhohrCF
i35PqD6q0Ha9DyVnFLE9jPDN4PcSENeAroOsukfn+/78tv9X9sSsDx/g6PTHLwgmCQLMLYd+nSFh
BumGVBBEKy2QQmO1O3no2eDeyC1W8gLVEtpWx9cYQniz/c82b93KWT+UpVmg9JxpaI77eeLkpYr+
cUMDHAO7H+cq5+JD8gjmI4bdS3q32vsDo5HPfAOnUTLeMXZ38h8qGlPi4uP9HCitIdAcp7NidFLB
JWx4vevW/DVKq2XHZNkTzzYmDHyrAOLsWuv3Ix7JBoZFvI+5PJZ3KsFSZ0vYeIkc4+DGBcDNHeds
gwbzuLVYaAQ6Gi5oAlg23545jvibiBowFkt88aUNZbqVRZHwIFR8FnQrupCzPWzi2pMGZ9XkVwQI
DBOh5rrqCqvjxDvsPspp9n91DWyPwYTuWZmZaeh8geA2rTiS1UfjizbSOntkpMIb3DGp2+B+h7t9
vIU/kdhKnpTO5pcM7Tso473lXEI+rddOuCj+6K24ap2yBFAkv7ZVh/0Dj9Wf650BuLyA/l7fWgew
zv96WQsCuYg5YV/OFa4nx5ZRFjDfRDIGr2Rp7x11jU+zImudCp6RgJf3DYraR1SYtqerkw+B6O+e
Q6ZsZFV3is2uA5Ic/ZojmQrlVTVnR6wT6NznjG/lDQxePTxbtIn65qql0I9XNeyAbEMoHGs8FQTo
4SeGDk29MMlIcaoYAW6kCHUTpZ62nfaF9Nv5ErqC8I0cYWp2KUrat0Y+V6iMxOXBw2zEQtYBA5Cg
Ld6KDwws6WBcyKdviZ14MEpoTUpwxW9KRBngVMc+YCE2JPawepKyhcjh5oc7VitaZuXGjZeUeu9m
loUQHZ1qJCdhjQ3vvKrR7YtP7RUJZs8sBo8O3nwG5SnFqyZGSAczzXMZ+XDjK5BSZxz0FMThq+c8
6KGozHg/30pGc43nnTU5Kh973RduIcNdjsThQzI8BlArf7K17saYc9tXYM8kSK/EySU8yPu2iUr4
iAqHK3VF7h4oJksz3Muv/FsJ7LAjwqGnQuSim4iH4bVPT4bFZkQIPG7ByO1ZBCNynLOtnr80Eb/W
yLg+L4oHxEJ+X6EK3LcRtRBDcKpHWzuM5A/w7nxvKvN7rmXB6nNCInsIqIZQXMX46esijXOLtJVx
UEcubQF1iZTQeVB9C1Yjq8tyV7fYGnyhrDsO7ggTvUIQprrqVVA/0APnNbH6C7b+dxtxpk45YVhw
yfQBayFL16oWxZ5Mo3HVwRAWoCNcdIuCEdaYf5hh53KMB6Rv4oK9O1c7h2z74qxLi99P/w1b29eO
sfiGH5wFWmfmZFUc1C0QP7TIBmAaQiuY8KRsxFIIenau3+8Lcd3P0CEFOqj3+wGnmS8BG/KVstex
KkcYtX40beoQDW+rciyfbyYYFCnhN1QNVX7s4XcOT0Xocs2Xj0obk0tE+XfJkV5Jvwngmx0QZxCi
09VRtCsbM9g3cEP8lafMfw79i0vjZnEMY6otU+zMWuN5ie4gGd+uKE8F94qghdW0W4z15kEiD2JO
SlDgk0vO4XXx43md5OfbD1UCitznxpDYLBDhXLAO1busyBLJx1VcGhwgVMrJ35u2XhGoHc3g80Eo
7bC2qO4aBZu4NsRq021UokxCHwCWtDzxic5DS0ouEKS2idnc3lVCyGErNkGpgyyo/06NH/Y+3n+6
KLjsBxSL51MNzCGUdgSoLLtUGPp1uKs3uyC7y3HBHli20XgddDafB+JoVm0LN1coCVu/Jm+9WSi0
b1Oxr/gN8v5fsz2uQksOqWUmLjxLi5xROQAfmpNckFqucIgr23a64pvzKYQ6NRcofLCQwuxcC9sg
IhCvUulHC0s0W/sTYnlhgmkvkrpPWvClpPZTOSL97aoXKxAbmFtWixbgKd6tPOkUtk07dSY3FIxe
IC4WCUbpTisPpwZPstg9sL2gEA/dAvd55+k+5M+29rEoTyH6zjRndR9eNIe9SHBwh2Pj1XSPP9WO
N1ujwrOxUCbMiwgshoDnErn/QCnwDnuiORFLXHX1zkZNeDZofdn7iE6MAlgi5K4bMWyQs6PiSWv/
PmYPV1mL+1au66dDLVtVMJ4rmCdwboBeCA+yQHFw0s9+xRR5U/YUVaQ47jamOa1wHfl0z17VKgoP
Ej499Cpbof2nbZOgi/LI9k7logh7ZNs0etg49LY9bMKdryu4VlgT4l9zYRPRe1brcbAZzpW89gP2
vki5rtd9ip3Bt/R4RyIsnwV5UW5MQjE1G2hiKZU+eAJRx/eEZjzlz/5U8GBFRVviKGYrlrStN2Oy
l5SVpi0nJC1yRbqpDl7MdJ49C/bUWEYFlv+c6wKqThidk8+409qJ7i23B292uMugiL6z/M6KzQWa
kQlxc0ZGd7Qwi/1C88YI9VFl5AaDtjOMVOEr/plB7gbCQsiiXdd5+6VdcHAMOl5DQzTaD+/TgR84
d+/YEYbcgvos1XamDx5QE7YWMF4PSY6LH+8JhHUVS6/wmD5pwSd/4eiov3qpl2K4m/8mlzzjvUq8
Z+B8dy4Bqv6pOrj+BQaSyFiJmvYm5vBKh8BYgHfkNCOMZFNYsEqQKeR9BA6Czkt15It5n7bqNO3/
2mZJBcZtKk0Itp3uTUmxJgxg99RHC5LrvFyp/lC0SCOJ7DjSbVe6ctVrIpOpUt5PVrqmpZS9QVL+
GoarszMN4KqDCR7LD3jRE1yOTY1CZZ3GHX+XnJtPWxXfdbo3l6D0QFNcFEVqvj5wvzo3FR3Qrk2F
sRdOeIpc8JUwCX34eMY2YHGkE60nyoWmWr7hTgoWJsa6Ni9duH40nGpEUrL00p9iXkBKnRmz8VCK
BY8t/hPsHDg7bDK92yJkUOEQev0eovIvNVf/TXg5H34RxFL1/hKV9/NY2vhV/cRekIE3e2rjEKis
xyvTVFeac1EQj+aP7W2vOht+WK1rb0BQdsdKtbku2ImWld8VY2lZQ81cN+3+owojZI3pj9RAhfvJ
DhCye/ym0QvjuZDMvgJhOPT5zPl9oCeLCbUDb+QreTJrD7ovaV0bcgYY3FdIhwDjrLRQWwUopZTo
QN9TdRXsfmkCJpCtfJ+t4IbqZsTxIqwWw0hQV7Qph/gCeSyAKOMWaJAqjuuR2+R2Uognc8x6+c6V
FAtPNaK5Zlvd6LpZR+daddSbkPaYLOmseSKy5zNBhyz+FdHh2wk2CONRBBJLxp8yoinu5YaEylU/
ROy/hcvtsqWEudbFP8PHEPnsNBMR8qgPSc9STjN9hZruGtVs8pM2yFDKQ0jeDjhYJMtAWZp6bgtO
Xgu8xtcdrUXcbni4PyEN4s5yRk1nAhZmyrhrfiFDSrxte1Y40WH+W6LeN12n2fyPUoeQ2zudfVC/
X6JweMOD78zBcvufBPMTm997LHsx7KMEJuKHLRT2VjqDVwNC5c+eGt1/V0481jGXB71XDBBTwNbl
tz+3xrbCCbHOzeLwASWHDFlptZh25DGows2QUfaEaPgg3gDbQ773Q0fGyl4V6hBAZY9FDPwRX18K
wzT7KmBwKHYjNcZdXqRRqMqbrhqxoN1OQ70/nIkhm2xtterWLk6qFxRwl9rut4nfIoLPurd8I3Qs
wkJuDEN0lNhaXB7eEdvjNZlHZKn9P9n9cKMeLhxkMrhU0q2u2nOFKuR2pFyC292NSFKR6Z2ZKQb/
fgAXm0+Z2oxH6lB+KyklBw86aXn1yVGIt/H/jJuW/qcRBoypqs4rbiX+iBnFsqKoLjIZQJljt0jG
Xs27o3Mi1L9cb7Q9btw3tNdF0GQXyFkr3Mx01RLdywKPKhO35PVDF1YfZczuWVJKSlD0E8pXMSFQ
NAW3ZKTCKJ1Wvk7jQ99j4DkjKA3e4OkeljQEQ6ae44iIcNKkFDm/OewiWtpjtrHEyUQIYB5pNCTE
wkbFsuFqnNQqNzoZdrFpSHdJCifo0AYuBGychE5AJuBUnsUUYn4feIRndzEj3p9kgyMi0hsNBN1b
Ciqxfxs13ERrs9ya0wZT6TY62zjegByCJ/7iesKAcR8h9InO6Qr8b/uryVs3ebiWXJb8cRZN+b21
KoDKJDpE4jfF4R4X/+LU9NjmKCZUNfHLO27uYnBHrlZRYKrp56ulkGdd2u/9dAitLU7CL2tqw92Q
Tz95xrRkos4NlY+6C3+DZfJ3lZuv3Mr+HW6gqmJ0tgredcYkgQiGb/BKHIV+VRUGnZxHLgcbPjaQ
Q6k/6l/ou5tWx0Bue3AnvIxPMjaNj/n9zPKfCpjlvLVRt8DKWIQXbOlUPJqhTxJwlRwgz2a++SnE
nh+D0Jj5B3Nor2CU8vsePxRqeU5DnSNzaluZFWKohSTuM39yYVNW2MkMDCNpZaNSC3vim9MqJvoc
KRV8wLPa4p1iYRzxAQY/uwiAtMtLCmmNIX5HusUTBCOIq0nproiwIjTlbH/goJUgtoqpjzv45XwO
MqY2AHlrNoSqnU8e1MrA3UhjsSa1IsXNISVB/EbwSmJS4fJ5TR42WW3iJc5R15Rz6a/DKeyGdQwN
avYa9B/QACYf1ys2hZjbtyqtTWmDLIyxFjIB3LcNmiNACQsGfmvfOSIyVZup3YpFZM3NwecL/upc
dMU4qmwBfa64mOMgy+MWm5yFj3XfONYBcq5GJJD3ugQy8wVWFECjGImFLr5sU5xOMtTMS6sohdNI
tFlYImYgWQQPhtHWBR2qSf+kCkGWuGBKdrfYYCvIOjvRx3cVt35DBSYREUEMEmlZyL4H//niNHGS
SszvmB7Mrlk3fqGrilsYTp9vabqn2H8OhKR1PiPaUQc2gx48M2+D18u0AFUIOEpnfjTIDDQuuvvp
ImOWlOVYv7JCnVLTa8d6SiW8kLgOQxzS/c2zx/N9qYWxAytOO+5hbSA3WfY0tjAlj8RipUboM4vQ
WdHFVuiVclsif8CN/7iMoFLq81bQeQmKZsnWFzP4gg2KO3NGdxnKN+Zi1fHw6YbXdrYQ2uAKGHsk
NwtTWvAMrIy/KQw/FRz6ldIJ0GvY3EYSTKEVoTQEtKlE+MpkWgU/YPPri9pxPsuNgXgc9DNBv0xZ
wTZxGUcbNRZMwxLMKpDFKi/ad16S7NxLeEKPcp58i51yx8ZBDM5L5bHGs+MVdniAbjvBRXgEAy9Y
7xF5n41ZyV1L68WhRMDaet4I1SqECLl3OAcwJOUGc1yL1Du3jcDSwZv0Wm+ps9FgCJu6BRQPm787
gDvZViGI6uL0epIj0fmsUvUIFSv+qBkJm1xzjDXJfA5fUkpiJvqzep+OreQcbxlp6/STyTOl5m+L
GsByDrwq/Sm/KC75pTnyyNhgZsksgxdTBc1+T21dEF8TkC+TprxGRnt35MuDxCWHhJyY6EcL/KV3
BRklly8pj4JeN4yWKY2ZeQbqjTdPyazBD3TZXtz8DGBuNwD9jUaKNvY987IbFcsVqaDOVIQaSWnG
THv3zxG4g6yM3e/mq9n62YpGD4/5R2Ix4u7th5DR+Rd6ynKUauU4PbFwHz8o8vL3nuQJrXUuK3U/
FG6ipsLcSqs4kUhgcPVKawOqtOtqEZLJFhoZzxNE/NqJmE9IyLw1Hg7DQMv+aL1FLcd/KoOj+PEP
CmOWIeSbsPaY6WmXJ9BcQk7glf8WRrpLo+Z+pJppDfWFtpnbGDCsZauek3SfgA2b6v07LObhvA19
2iTqGKOiWdh0G1vGEZXVBcx/roU8QWyozR5GY+8I8O6il/37CMokVcgMU4sArOfQ/Y0FSieIuQWH
PWRs9sOeikPOrxAfE8VN0WDaexyK9AFfl6DCHKo303zVuNI3Z8ofuH1ZiGol9+tOXIv+sPPBRPNe
NbKiqd1mdhkp1eHHQ2H6Ve2hm6HVIsRyW04DBcpIyYJXv1Lo5kRMnKxiuf6lXi8+T9+bv2rYA36V
bBNfZGD1yhRzpPAEIl9ngiklXUlm0kUlgKZpLPg/AEjS2Mr7za0P+A/18G6vy4Lt0UOfbSKTAU15
rvrVTJpYkPpgI9MmRLRO80oTD6Ylt2x71mhXTRJ+tfSk2flGk53xQT9eAsSvdFDjmLUVkg/sKGen
4OihiMy5X3cpA6fEucX4epE+zOxRB7eyoX6B7XiisS+J2fx+EExJIhpAuznykwOJxQ7gA0+gEtPT
MOZ5yWZQozpcZ+3rya7DwtNIDgpOTOI9pFhMO9gTcF/tu2z5BhFrzWMc7EWmfu1CCnSIVfOTuZu4
UMqBEqY8n+rVKpt2pACv6x6D2rmoGnC4c/R282C96wWKt2Y2JTeNauFHZ6BoRmJoMj0Don2MlE0c
qw7NRSKSeMRk4XyTpfczpW4eup2jd50kyMjXAiAtGzZzjevE3dRvWFw6/6tYjVf7+jKjKF4skGQH
AJpiDX5jRSDdGhkfhlhRQp0NapmCeg+7iHcvADWaPcPpQK5bMHGDYZ4unRB7YglyU0X/HrbIxY4I
2p98RkWsPjBlQkyP+/vKUZ1SQuqIpNf/q38I/HfrL7oZhYuQMtpdaOr27hFtrGD26P9UjRgLNHSz
kpfFq/Bv5f2+u9GiAXceBpEsQrsKsky92slBK5amr3I8oJi2hrwBlmh0AZdwOT8vlCji7Yi1TBuY
e/nlZneJva7Bc6Icrf6cOt9vg/Yy/uoE7wI5mzpsblzqDAG6PQUq64maaI/Btakq5s5WnpYrg5Xl
6OsKAs2h6xtzbO3mqZjc9lADpNZha0Gjt9tIEBNddMM4/vYHLvIxwLAg6A3gvM8ik2Az+cJXMEA3
9U7QQHM4enmGwGUvsmDfOO2dLk2QDqaOX/XYdWta13RN4e7/mWBxRkhsLWYcYnSVIpRDWIr8IyJ/
Go7z5P14SXRphu4hUp4Pj+V4cQ+gptNLuIJbpWDl1XmE6GMrZozF5T+tzoHAUUpKsaLYqJ5qUN6k
q2haluhnhnwwxSkhrHO4LMILIsGXgOLvcIsuLMwtSHEfnhUgdg92b/iVh0wl2fvV+YI7uuMSQ0VM
peRt/xYZjsR7rtH6r2lu3Id+DQkE53YJm1r8YIw8bC5lDpdyAUKHzCq4m3xzcZoK+PJSy1qf8Ddp
C9TiweuWpQbOEwvINLq3mVjE11iQhe3EGJUnyxawESijPsIsVpjykPwOLuZ80mO3XrNwBvKsKFME
gUFx472OTtADOcP3rvBANauUj5E2mgpN10L1zl+zirgOLFOAdxRzK1CfJyI+fnPEFD7N1S/UInSc
bvpUGLDUrCFNJhEuYanuR32DZSG9Jr0zJv7HQTR+izxEF9J7YFvrsMCdlZ/dQZemGjEpc6FcFJSZ
MMB9vpmG3kvkh1BcEMbDDmy27cuIc0hdpc3lUeMcugZ+3KXK7syPPV0fKB1ClZRc4aYuJgHq7cBX
h4JVg8LejHXgoUsBnXwMksi9g8rhb31oNlQfLtM+ChYj0hC5D1V2vLL9pPR92N2X4AaMpCvhOSdf
dhYvOGhnKU0/zHpkOtNvtK2AxhM2ZD50RjVHsSh+yC/Zry1P7UCmoMffyhp1JgG8SV26HUFKr1Ku
Y8dLz5xWtoGlAfYx6NL9w+NRbhMrI4Vz9Be8GCxKc26/8H4KxYjp/SXLsG+maH24iNINtrz5o4By
NGLNSfm/GfTZbuZjNtCSZKL2gnwjC+rvwuH+KHfbXTi4rd3qZ44PD7nPo6wXzjt+OUI12Pth7BSa
PKH7TznE8Ik0Hfm8CFw1eDnWzTynKMVZNWcDwx93nsyM0+oQR0GPCKHclUoySnQkJ7tSLjbVgFhH
zu5w045YzGqcgAhDWv3mywk7y75rlIJYa6e3HaWfWfDBrHrbrJydgeqEQ/e+z2eSKtz7UrgDw4Yq
98tHZ73YuLYMGQjMsmmQu04OmNoZJgkJjeSeAL7cWE87Lwm8dwU51dXxmcJriHrYzXyH2aM+ZojT
cYFXCy1CfDBzjJ8fe/xJe9xiLOTAkAClQy933g3Myg1+HcPrH2H0h454Ss6tl6dD53g1H3ECO1Gs
7UPex6IYB8GOkbYzFHkK+5t9+tFMusudpncQobjte0gZzgrhS3AIUs105o26EwvNs4xgez9URdpQ
yfDqpFDikpfaM3oH+rGeGAFGkbBWObUz5sK6h9cP7Eri1/Iuy4uqz0OepJ/U2UxjPYFRgptlQQJq
BiFlz2hJyxfVbd37FPfn8FcZPcqUeqbECZD46ApxFgMOLXphY6JWlehj8Gv8EcDPkmi1GC1V6adG
EK8QX5yYZWkKqWzNGm6O0qjP5IWL9jcra1iPDpD0FtR0EWv73LmLDiEZpwMjMT6Xn+Tce3gCns0R
FCYBQBfNXWlzRC1yW/c0ZOj86uGovqtykMk7e2S8ovANluNyzyuUr+SWjcf0IkmqadICy1EtTUD3
7NxzsLr+Ckz/VdZmi2vL1FxAY4qaZYHxsvbMGDFP9rU+3AxHQx91enBV77tvFFQxiyddE2DrDbcm
IN66VgzuyHmETCWnHvPL9rFkxqvNbMzQpvZLzuZjagnH+9R9JzH6IxChaWj0Pu/T0XNOj0K1e4SC
aBlo1gCkxhN/hpO85dwo/JOBnCGCdyy8b2i62qT6iwatM84Io5Y7Y+thOGttrMEVBxknOi6HeQU8
4zTmFkAaJLbb3ZAw7XSx3DMiiQhCzM5pKljAGmFOwoOh1t758p5LnWRxQ07vDi5rp6bIWNgqDhGc
tmVhU/PFnZkxoV22G3UQkR7IMLuHdSyffv6fJwhWAohf1WrWZ2XB+wasXA5+63xPPdP2MydBmK7A
4nbasrPPcOkfxJHrWLuA7jxX7vuhgniTNn3Qt2ie7IuLbG/hJOq8f2KHi0Z51+K5Zwsapn+grZR+
3NNFZsb6iZLkNLltIOYmwSYodJlRjW79pWz6Nbe+ynRzfEP4O0471VvAiccbxFRSh38e/AqUsyhS
j69zHtsCQRZ6xtioRNOPzeApb1OeLJvBa5C5Yu1NRu148RaSTxxInsgxhSdJMmhrZp4ZnGkU1GmT
/lBHrCLxRNKrzlhoxhFGFrHLpns4fVbRQY7gB4H54diNjpzxybZDJ1n6qUTUmXnhtNdQUP/Hju6t
DjBojoR5E/eQp18kAF6wGE8AueSlSw5cD1EpdzM4Aj5tfAsnIxcMC17U7s4o4W6ija7FkmRdkcy8
BlC8oYxwzvn9xuv715cX/FtQnEpGDBksTUre4fvfWAh1Hw/4ZO2V6J+pT0VMnGIULnX535hRCRwS
G+wCDl86RtDherrig/HKhMCYlDZnmdKLUyOreC+t69Eg/RoWDjJeEHrjgKqJuzlDwwjGB+1gH23e
RE7dZLpsvHPybMaN/WvES84/qoVNFuHqf0JzbyQQ4HtgvvgHzFoT+/iS55/s813oHd7vUkKgR9KG
i1Qc5Aq2HPInbdLAViH15tQG7cV9uvQ/zQSUCHi7q3J51g7gyFsJP0ZD7LDNgq8+njMdbPetWFhu
HCH2PJwOXXV3+L+s9eqWjaKdvrxKEMp92JAFwN5FUsMGK0WoPV99qIWKwAebSrFC18vgKpo6lbu+
1CDiLVG1b+gQwnX5Frz+HdLSajqUdA26/ejoyNVehThocSySWCd6vJdmfpT5JwTBAHtz9lPZHaya
n29dLWIBegLw5i9dcmUMwGwerNsjAm1vIFm5O/HFZw5m4wYATdBTS1UM0B3mAlLd1wCFYiRkg3et
5N5kK1/am0OzuGoRe8H5k+FfhHCOcAH7Uklut7coqez6L9p9HYe/Mr192rfqxeKE0wrKph6CjjV0
3YaLGKAz5K/HwXl68dDPpDC0V63x3yJ3lSoj4Q06XnYKso/fM0n/QDDZkEsvAXll8w8/Uu4L1ayr
pDo4vivMtglLbHh4/8iQiEf19dsYUSV0l6g+9hkWksWl9+GebuYKNiBNSY2kQC6SMStmBY5VHlvK
utqUTJ7phw/bowIRT3dJNLsy2QhJVvbzA3Ao/YPf8AnQul7jts0BNM19JZYfeGdLnm9HL2QOR0lz
0odVKlc/3UlCb951SfG1+unAB6xszNK51QbqlU+cv3LMO2dQ0DdEsoijJo1Q3HjoML5HBKjewpdg
WEksa83UzGhHQXR3quGvfQzrZ+50oWMM0GoLVKzRBM02khJHzH050J4rin0yPPlG0p4vX6817UBw
/Zu+CJ3mmcK3WsJKl02Wrf4KTWXMQJNDrvJn7ZEj1RuUQv9xw82ukuGLWlE7UlqVXnKWa0S0FBNj
PQgnhsXKSsEjwpbOgBe2VxM537tOlkD+0UVhZ2TFRDPbf6/pdwSDpPwRQC3va3I+cxreRa2W5i2e
h7mBOZ2RXV0GnCAYiOIi5/gmlW8WynwVScrdkX4othf8e1GkkD+0d0ewg8Qbu5VgUVkIDu81/wXn
TfkUU/L72/KUMB5bTfd/vTI2bhnYH4vSCE9ax6tLx19dxxNO+KRuTfRdqKQ8OnTYbiUCpF2vhkjB
M7XI1G1atTltMOo0FX2bIJM9ljFR2tyWRrkSkNRVKv8h3VUcqdAT8aDbCefIrbzjCJqIhFIxMylA
9MSl265lKLbjjBaOd0zDGL5vRXKUH8ADYeqbF5wVJe+YDF5OZ6E09JCajQ4DY9nW23WvFkRvbCTU
w9ejMNYMcbhdVEKkWi8wmaXKXPoJ2nJSZdd1/0DwInT9dR2zyJJp+2o4Iz1oXOxIuhc2Xr0KzGA7
YaCcvBGvz8AqPNyXMrWeDrai04GRs5dcRJjWIOFSr0xwBjV+X/45Oa+ZZs5dckak37jh4E604M6x
4DUYVwCuuiDSoyLeLTKcrbcoAghvvnOMxFFhVew7xe1eHluvUDOL+XyXZxV1iacBaPNcEzSSpEPn
/RlP6o2Mrn2nrxdkin+qaO7qIfvl7g2n3uD2pETo1wBEQlhKZqA3u4FGZnuc4OKwVcZ6J/D6Z4U7
x2hP8Iqr/NuPigCbBozCWO/fOLekxFmxom7sb7Mvy+R0SAPIMDdJ8Aftb8iCQ9KuokX9JcqmOqvR
c4Ek/RKr5mOBEk48UulXsTk6jwOS3TajWXn1EVbgA7zLUOA1EyzMGTm8L6J/EUIDWEvIlczjdabS
y4K14mfYVh0rETBdnGuuzruCrsTbhivud5hc0MlldmSB7FIdGm/z08yeWoMeCcNqjy5hyCiE4ZoN
V78R67+Umhg8MCPKu7E9UQM3v+rQQ3iwAHtTGmwSC76uejPwHiTvKIxHP/76otxuZ7ZvP271da8/
XpwNvG+PtdLNBa8eA8dhL2V3Vdq3dHnyRjv62Pj02S39Jgsr/jTBuGcMAQmcESgiv37z34imE2BN
lE5TlSJJTNUIHO4K4G8992AX8dRCVfVwoOlJ7EGQSMPgxrW6PldPwPo8jW2YfenT7NU9PQpG0O8M
XEogBwdI+SC0KD7zjRk+YJMnB1esZlNNGoOF7PkBLVn6boNQhyc+oh5O71/F8w8acLLncCEAwuN9
ZC2IR+DTCbYY2FZMyL28bbxJnlkTgSxtaVARr8IGpCZ3pnLblXSuhfrGjnDyRea4DmNPbDE42kmi
52g5chVTV9Vg9J5y4h89dtEsgAaA4iGnodKh5Y5UcZx/KlAthdGLbqulPRPL+ILUxvqWC3LQqgGL
zWd79myWsaJo7evayklYG+waNRjYRy8nvMF85hHjS48SDjEwYNLcuztzFimJ7gi3D2tmPQvWnDdf
MtNgzDKudV56F7fxyMB+OmziM1k/80oh8wsHsSJiG0CnlOaDmLKA8+9mbB1ZOSpDN5+O7c+d98kL
rfTLjEI2GU/2M/fKeDag5k7gMspknP1x4aWppNppz0POdSjPtRPZcL++F2k/9zTt8EB/FaxuSjPl
6Vg1YyF5uLisdntS/9NJkC59CTJgJJH2/eUu+AcXEdYf7IgRC1vd2aNSkwxEWCcnX3qeoyQ2VvEG
VNg6YfEIZ77s3nsaKMsQ1EMfo4zH8sLc/raygiZYvOY/di1DycTATOUcvWWG4vIJmpueh8fpM1LV
oxUsXhLUeeNgDhOWNO+SkL4uWmu2B9T0F2HBtUORBlldOesgqyEnHUAkn6jPOub8iOouSO68GjZ8
qTjGJOcwyt7kG+JHqI3cOyv/1hZtIxM3VHpdYpxMRfufo1jJIzhcvfyQkW82+nzSZ2oYOMBq748k
4SMQm4qYfP5tLIN88YijPzuBFiMYZOAqTyi67sA4nsiptGzbjUk5PdPIwNtYu6IWTDxTTcK/ALi6
gw+GPT9zbw7L9cPp1BLRt0zTn/G3ZjbHyeLSDnwqA/xHWj51eWjO2buoyqoj7hhroqQu6us5Mqal
fyEJmAvG38kshwUaxltZ8zXYKJ8BQL5nv8HsptSMoDsfUxMAos4DkvRZXzr8HyFZpOOhIqORpKXO
3AIovbn0KQ4feoW/Su8YiCKnhh6qi7ipdnGlP/MFjagsDxX7UvBFUoEwqHAG9kR8dEGC4LID9wPt
9e5+c/tTrEj5iGW/guxbu9vaul7zeEYIy3xgNgMTfT9VQRZ7WGg45fq2M/6pgOmUFFGXre6y/K3X
PyV0dicmCZTXtuA7AKyIMDOqPc/Ji7ocgavHvt7hqBC+TrjVdxAa6/m4/tKsyL2bTEl/EXAW+RhM
zxYScQtXI36C8nmc7ahTHS9hK/93slTvnM1AB6QxEMAbtFa/YEOoeONfgDIwh5HMnKSMwuX7J5Kt
r14DjkmQlUKdGsbV9ARHMSYU8jvwclJNTz8s1H6awIltuejX/jHYpexmXg0LY1nRfEwBhkaL4Jit
ctTxTBe10CywOVHSAI639bmsvwLcrOMrzK8EG8K+QTgYtF3btIvLi9fXl6EmkdGc/s3upeKod4LH
GzQZxrmGIHbdufvHQrH4ISlRq3wcii8fwMDyURPIFHpo85//dD9SZ1mVzY5KHYmvp5vcSrjD47XW
1mABBwkwDPDuPwYp2WSSOWx7BTdedyUoOZiNcS3tsQOwykra5UIL5tPu9zaxHpJkuD4R8kzGhGNv
Ff6XYEpgv1N5SCp1djHzh5SoTmQlfVVGLuxz8VKppHcrcqAl1Iq/TMExFCIy3dVQCvPB1X0XMIG4
cX7DesJsajfmIyCoyVawtxpGc8K182i6SYEj4TwuHDD2INIKz99XOdd2jHcpGVgyEqwe9NYKcLHc
8n0baQLI61/cxg6/LYaAGRlS6Byp2U4OsovH29BZsP5eBY1jyj3uYELIK2/UJxoJY+1aLYqwaAk+
OD4we1Qz9dEGYjuAT+X0tW7hHVd4uqZzE6ILFnWFhaSSdm+BL1v505YUFKAnN9NAzcTuTPJLzCgF
KEhBX+PLyEtyQh4QPwki+2f7RezmGmk27FOjRaW8jhPDCJOrD+rw9+kEFfvGtN18c/i5jxWVXivf
f5u9A1AiO+oaEpRTQ1ofhHFnsFFFTlhYzfOI6Ctn/RWBdhWgvl/ggjKiVARC0JoeOzpkdZHICNzE
SPa5i8iNi/jTx9lQLsOW8NAtaJPHn3DwpHhLjZy0CVv3WDDV8/fXs4+vwEkgEa1i4zrDnd9paK7C
UXVBMWIkdpaWuTj9KSmmzJ6RuZugxJFq42sXfCYIoktzq22HRTp0U+xySPsOHa3997wXfj5N+9mb
0gzrhgOEXDBcH0kKUPOc6qA+JE5B8zx/Fhw3RQIuzfKGOPyfuRV/Lx5NQONLJnjRXffxhoIIVlFT
bDDdA8pyLJnLADP2iuLArdygQjjIrg5Wu4ew6SKi9mHh30pTVioaDCN1GuOFPcdbfmpvN47IWJsO
6bK1gqwXGLBcVJXEt+3m0SQFvL9McebJHM4AGNMTMe4ZBFs7KgeafQG25Egp76zu6rrNVznywZXW
1fluEiMNtwFBjPh1rGlf5vacJco8ZkTjV+aCWh8YGXGs4XYlQ6YfoXU+QyUmX6FbMYEbu3yyEaZ7
BL1ehPIyI8lwT/wzaRyNCc9ZJXNGB93nhyQtmoslTQydStROE0EJTPtthSKB9900OGMgZW22Aetr
vTr3e4TSzC1NPdh6bhEP1t7NmeNeG8scK5ftPa8RUI/CR9npmMuxyujM5nEu/rztn/6SIofQsHl1
24xhuwlg3SRiJ6esP4KIjEZvCIFsxvl3H91Unb6eU4WSE58cyaJephase84bE5I3/6zuL4KA995u
rbL1f4jsxHw1m+Qf2UOKH6JA+07szpBbKMyCJpRB+PClQ60IOyl6sXvTfKW/P34ncNPbOvapN8yV
BfWR/v9z2a/ENyMQ7ILzJ6YC6oTbLZ0zijof2srUiHErr6WsE3ssF5CiW4s8LI2vRSlNx+MI9Vif
6hMylj7rRnUlvcrvg4xtNyIuITTxByvqvHhjb0HCMA+KdwW4gKUBecOv3JR7eI8gFYoP+q/SucgX
UkDaOBtlf0g79YWbvWD/tvlMwdhT0CStx1nvXTThUZ7r8j7IWF7PtVNPrI2Gt4wECIYjgB6GdNQl
8oX4+JPIjATpOtj5XNKYnlSmjnRAdaoWMhYQ7IhsJ2wToebqwXBJfMuh5uw4Fyaez1CM313SeIHA
20WZzAIwRKUL6Iz4gq/8tlZjeANVlZZ0diXX2+I2/I7QWl8+8myW0bBjrAd3LcMDTVQd+j1CR/sI
XLDJxektHVuFW7Pn5NwzOMgIWloxOqx5ESLlpEBT9V81bBnlhEJiRYgFFS46jjGwFo9hHXRJbW/k
bFCF3Ykvlk2gWD64VQIVO0AgcblEDVyJO/ZSkpy6hFo60wjsa59UrgLckkn6N5FLzKBBVc+EFiBj
ggN4a5Z/pz/4RsIVmunxSS78JPTZBtbOuqV2szfXkFao4dEWSo0TvKZfpN78haLXcSkc47Emd/l1
gq7cW0Krh0mur4IheUIsPO0g2BIWJuigGrCbsyfzEX9Gr22iPJg2f4F4ERVhDTJBYfbrSn/vB9yx
7nQ7nkAAgvvXyA2nne6+jY6FEK4RWUd9h+5LtIIw1BiKG9jl6Z1kR25AJ4fvc1NtzofFqS+S3p8j
14t45+J4KoJgJ2ErphzSclMMxdT2jE7OCkKScY3K3Zv5ktuyOQuF+2p5ucV/k4v+AVHsCasHqOny
eANs4U2hgR6stHvFVwjMy6sQYdmncJPvyavUdq7KmcVG5i5hWjXOg3jX73SxnSlRagl52tEgImGZ
5gtdtJc0G8fUuJCTyur4flIx/NtjP6mEUgSphLNV6XSoOd+I5mTIgVwcXAPZFifF6rvbPvhNjiZM
BjBfhCAvVyUZ+RymramZxWHwOwoGUkRk2bmcMMZZGmxhXUtrA/CNO9Oy7zgPbxzlQmSXaV+Y6Fgi
AXe/2j5WeSoJQJKN6JkdO0KQ4jFzLSuDNDtXwfvQa9VB0sljgmxIzqZVMgWkxrLdSlHAVHx4U6er
bPgJDqYHxyr3YsRacAYnETMvS1Y2uqgQC/00ToXf+EuF9xNlbGAh6+zDRLbCPQokkYIsx/Lsr7lU
2T4yPnXr3tQyOEeA3erwCbxC4mqSdrdhhfd8zhzpPI2M9sSU8LaZ5wnclw3Ig/krIj8pM0gMrMW0
zMv5jfrdTRZFymDAyXbsNM2uDWJazSWhdSHvygl6BtOq8azyIE8inOdO6yVdD9L9ZHY2PiLn3jMX
pdbsfZRFdTHbaEO8RPvwrr0HF8wIqvqS4gSLeXfO+mIi6Oomidwvc4fli+mD+blddEJg7SlfCjpl
LNB0i8EgByPK0IUfHs9hP54fE3O66TeA5wYHUZ/h+kXU+Uqa7EdH6GzlKdsLqMBYmFs6iY7iuQVx
NFywgCCyDt43y/GoSr1VJ+WXxxOD2ODfBD+maxI7GhOmiJUtVTvM90HFuoUfZXTaMAIseX9lCutJ
L3P29/gxGu8RM4oEuMe8jnz3KK18UtC1jVO2rdSFkJ0jV9/s68Kn006FxiMLqk2C4xM+/K74QYms
4/LPRDcOjvx4emDJspHnulN6ss5SDKSUloDIZjEgrKnHsX6K6CgO1V4ypTojZfgGOx4XR/oVHa00
K8xQFMY/8ELZEjgVUg3X9uyYK6ySvwn+MEPrmy0bg8Yy5Axybvd6DcudaD6UIl8m5u4ZjDt5j2+y
MGVql7boAmK8uIYNiaoFelHNsK/6s0DuIduIsSKzcw76tPmtp42azbCYVX65NsgT43Ql0R2w1Qv6
hmx8fovSzJi9CmRvoLuxGUtrnurUjMgFoRxneoeUnmOYqxlLSB/E1ePrnlf5928sUFLLx2uCbyIB
04bc/aQNLUmQX9F7cmDhH1YUCJ/G708pHzmcLdmZpjSyaVfSgbGOi6npZOyPBV5+u04+fEb9Mtfv
nsKCzdUOkWfRA5Fznnv5bkDCgY4CPwEZyAiZCiTqeIOigkH8FOlAY9NEYYMlbKggMNdeG2FihUuq
uCcpjPz7TqAFhQSAQuHIoy9uE110NAMC5E5didlMvSnGWvmRSLS+UfGLmVrSySvPtXQLpZYvSjbS
3be5czZBjZx3XzyLTk6G4DntOjyJy+B9YaqsL5Ta+FDocx1hyllppF6v9VRDG8e9o3G/mUeCJNMw
Y4j3hwYGV+92335QImd16nuQG12ZRO5ocW8HI6flw493qLC8sTfTHn+9GuRzvYNAIM2pySzQVZmG
xskOQIYMdUWbAZEnXQzpSxC0VUV8fxYMHN84Ntp57xGqhH81mu1RTq8sGE8pdxw+ZPGxSF9P40E7
pKvpCx2Wxj9uawCXOwOE2Q0eza/8RIdosbXqIoFG+JPFyjm75rZh8zJSw9HMQLsxbenf2MxjlfiD
sRrcAoNTB4nf3gNT2KvwlJKbBJLq2unqd81a60yU4C+/y6V4loQ4bGBCPjikY47iyBEQE1O2jUza
WcbwduKnj0OZl8rSXrB1LsmKCS08mQ3dhH39EVCvgklNzAmx0n4B8/RyF04rNz94JoQKdpYeHHXq
FPT38JRnCSrcQ1+bAsfx7mVwXsezLKkl6nbQiaXkjxKt2n50PP6nBQvxcw5f87RBWrFXsPQj2pmq
cWQCE43qmYluLjz67bteU/d+4Z2WXl6jPAwX0NbC5uSvNfgwU6TR9MMgfDaO5bUMSYLJdcE3H35q
s0MvXoKPDaK5iinPoQJkZUO6G6eVCcLxkszuGFiI3stzsZr+UgC4vV1bj0gniWRPAhaUcyI195yQ
7PgetJrlPv/8d2OP29q7DSXvTlkwwDo6Xwaw/KSpwDXTkrcLZb2JrtzrRFMAmxSU04rBWqZEAwPs
aWXaT924agOh/fyiyGs6uxRaUBwbOS6ZMudJmkmqgzX1LGP0QEHJBlrZHoo2D4z+5QjaPF7+6JAx
rDcsARM0L4WllQx7EdTn08/ymelGjhRzRncKU+7v8+xVl9THWl+i1Ml1ZLVwlpiSY7jm/iHh7jNE
apcfcUQEXMiQYghFcyHbtVSS4QMVF6nr12XCUmMoLwzL6IHei9sFJcSCRTRi0bcrDFmnq84KpIC7
9y/T556OEBgHw/Xs1GCSi38Wqz0zGuBKGidHedHW1crKhWkeq+YdMtGAJD7uwAcSJfFFQmXr05rC
svzVvbMJZjGM9rNufmo2a6vm6W8m9qUOuQTykTVoENwzJCJgCqx+RUz2/0A2c8bqjnPm5T8m09Oz
Zq7xUxPDDSIq79MdwYA8wS3QmBu40ayLP607NIp8uJAumDixtCCnfFEbOzW089gKd2t6D7Oqx1CZ
EeZc0qU2mSHrUx/mHTjcPGVYO4e+qr6PO0twfxoECfEfi9ediUL3BaWq69VlzJJbKmAmwlA4ZUh6
nPL/ewL3Ma9VGYalpRE1EsWUpkSSPNY3fUrPNGPekixOxTfjf0f9uJO7vTdaEj/Lfc5xAVZj3l28
Y3J83FZFWlfepEbsgxsLBa1nMqnyjUhtY44OAK/iGAXhQIYnd3mbsStvSuk8rp5iX0e8f/SxZ516
WtGjhJtkXK30syV2nmJejYU96QzJ7ZtcuMULgntyz0aSSLBCnN7gCwyYp0MJM9ng6nwxFX3RGHTQ
bQf+I4Sw8IzbPWjniUgs4x5ZZmdVJySTA57n2TtRuyIZq5CxRqweUq1GeBv0bk+IvJNesKCpZ3ND
ZwREccpwdWn7Qf8ndptAcamCnQz3+b/Nl9qZ3Oga4BvAXr+e9qivC4dAGTJRPcBbA70guY0o5oyF
JA/rW//VU8nbScMC+Z8HwlaoxcU5xVgewZsOQQreCPCbkMJ6kLLDRYS8qGggCcQXdliVRHpm/LWz
jjwtoW4GXbgHSZ1zKna0XyaMFFA6AvHWjgcg4FuoBTXBAH20aUlxr82rj+683WDIRj2vNbiGKAGd
G2A5qJ/N1NCMOTNGAS17UavrcX/qEKPatmbQw6oMLCJPNL3RO2K3jjD2bbtdM++Ung//R1yQAtlh
UEUwCPMjLXu19xbGV6C/3RuDjvxEs/AJneMj+86/GVUMDMzTxH27p+MzL32NAcKTCMjSORvXiDgF
yMzeN+FGbe3FMs61DkarlJaZVrO8+a+UjEEd1i58jgpvOt0aCYVeUnxPmtOj9Pub1ooue7s5qn3r
FojvU10jJ5/lqgttAN0VYiNyVdd3l08qSjBYUhfRGfXz6V0t1CrJNbeEDkQ+OnxZqLs805fZ+XQ/
nJcbH68dAemNArlNK+9JlNUwcyn4u4YM1XGoTGeGpIShlx+IG2VcKMBEp5N1f+xpctBjQ+oCAP4V
CP+YZ4XxxdPY16JiqQoe6JlKEsiuE6DSUYJxDoUbk2N84fsX9OFzQQu7XW/n8zBkGRKv2K6uLngp
hwfxyEwe6iPAxBBIX2KMQsyiPoywiKtXN6CDqaZpYTGjpEc43iVFeVgQYAsEJ+7X1xBRVvHY0Awh
SFAmouoi6nO6w/qQuJRAM52d9eUtv176XBTvcMUaRX+45cE2Ci4n/OlPnpandZYVrvoDrDyPBlbZ
QwOrTYrUefqwuJI1FxXyrPXz7yU2XTBlaiujmRUleAr/eqw+sowFaD2WhQi8e6vHQjWIdBJN3cFc
z2T482epKTNVa1O6VkE1R06ndsaNKVFMAEtSb1UDiufzB9nQDPsdbWMz1+nBbcax/dcQgbqZ+pEo
0mMF/yHEkfzb8UdOF2gJH2mO2Kxg77ObCelFUBxBM38KxKJiNv2DeZPBLqpCf18aRb/fHUAkPTIq
+mt9C5jXXZowO1jR0O/yipIMZ1jtbhJwnZOzlxKAeErOH3Nh6mhTIbjEr8xfxw3fHvZfy9jCgG7I
Hh46nZ0ShgIcII1ixfngOj2piLVqU6Ke6H/fIKWbcdahQnwnKgsw5aLkSiEuLZSdalPaCnh6bnZf
LrJqZOAqwJ2tq1bwXrXGq/8nyGMLGAR2WQ2ay/CyuckPZMwQkwbtoLmzAoym9xGvb1Mo6ldhf7yr
dcwVIGHXNdOpv4TzY4QzX5e83CLqGv9xN0/JocUWaLFmdH2GtkBfXVYRhrk3OlSC5iN2tlyPXPwh
ZWzALuV5e0b+4q5Vz+TsNbmtOZ4sb2b9FwPQm0/bMfk0FYwEm+pIiprdcmO231sDWP7NNAJY8t/8
BjJXmiHghrDofQcEjTvXhajQU2fXylsY0tK/E1keek6h/zkghO9K+d71bEi1xyZH34+VcSnVVz0r
YhXdwcFmnYcKeSKa+J8HvfYbPSql/XOUKgxnPLavJ5mvZgWHG1QEz9lddTotxZf9PTCm6+YE20hN
LF2ua8SjadTmdxvR1qzxIeY/lUNPt5ZgtKJ8/Vw+0rCN40KAHM24JR4kqKVFSq+txX5nDHEID1zl
qbDRgvei+hPTRM3bq8aAg7YrVJKWtz7AYAGY3h4ouTFOOzVN7dSzYnzJDGxWpmJyNWJbUPNovvTS
3z5jfRFo7vKpXUBKSYCFaecmmiF2jdZxUX5FinQ92AtnuMyattlxXNIsmMg053QNWGzOlIcfJy/7
ezSEFvdq9wrDOdTtjxAMQhUqriAbGDA7uMGvmOchEHZ1wj+LLcLaGxz2PBBdtQ/fIyGmS/e0JUxz
0FBfdXA6Q+uTz0eRVGxnhUarkE9SzIdKiQvq3Mfq7TdRVp7/YiQihBSf65oF9J2KewqdnMg6temP
ZZpoOygSiHtcg7dpktxhuQH1Az9g+1Iw7cW1BzADmkbU12RtWu70Zlby/aJL1lkFo3DqTCpbejix
ux/3kVGYEjLGJluUV+izn9sYkpQzpH6Q7AnJ8hCFiuZqfXLH6oSWnRyK1NWGH2350fzi8/S5A/Fr
MtsDQZo1YroxLLYOxQf9lSmZg85mQgHTGTYQVmoUFQohMI5PbgaB1GQqSwJYmitdCCSEeandjlQz
M7ryiirmX8xFwmUNsvVDcalzhA4qd7pdXMAM4dq8Zo2c12rMcwr3pJyXsjDjfX8eRZP+cb3Noadw
y0LETF2vpxxkqUjCvYGyvO7eEKY2mTeeQW2dU4mXkRMW6VlYJmodG8b7XUSl5mU7I4FBjjqkIEfJ
sHBoW8kW9QYgPxUVMBTwZIHQaIq9rY2LtByjjjzvzy2hh11leiK0ud3P6dUGp/LZxg39vW3NZZ+e
B5PilOnPII7980y5WLuA+XB9m/w4AosCTomPHUgjqfss891as+EY9mw98PGReenq2+uPis5+XlBw
L+dTwy8qOCyWyNQ1gGu8iIffJ/lxLgllwYEo6xzyXjgAnpq+r+fb6gwgi9GK3GQDEoQyhx4Jz8ly
HcBN3iCS8IL51p0pA7vdxQ6ZCStrZRVq2RRFKvnuX0oWMiFs8e1NO25uT53gsMh1w6OPOeBxkO4j
bsRgag3CRg2nVjLHBt4gqTUsfbt0p1G7OM/c+jVhy8C8q/hcbSalkCehhAJDu3fkuV7sahZzD/xN
MsjhxVuycA4fovv4e2qb7tj6DR66K9Eibab+Og0xY4Hg/iGQSS6oXVDeYMoBlizR4UifkUZN5qA/
k3YjwUVgRRI0vLWvfeejpOTfvxgSXb2VYGuC9/VKlHqOFYudiHUrGlCMpJoXh2FZx0lrpbFyA15N
jEa1c9KhVPKK9LaKYf04dJE5g19H3GCxLmdwmr2zGjGLfq/xZoPUXTy2W0c8HBo6+2Rti/EHN78k
CYvrUrOAlKzwi0P5ke6tSZJdGzYluLPvLo7zSz1TrTv0Z53Q9qhXlgRdc3AH87QDuicy7u3Ypzha
KTwGiz6nkfhuPu5thZ8WZVmtnAoldASYxnRdyLblJgSmRNwRhhfj/r4r5QDCEkRrUuJGIFtcJmXZ
cqyf6CYYhpbhmLIzsbY2YJ+GlaxRnJJ2u4lU8STWPp3byej8KGB912xX3IqvYOrh/Mm16bzWX5TG
SL0BcxRK+V73T6OQwCgj0odxb0o5VrQ0ohfuL08orNHSfYExIeEDJvYTz8mHAw4GlCxaR15pErD0
mgcF2O2z1xSVxRGJNy8U3iWopjOfYXFB/soeht4ofvCiT7a7r46OLzBkp1fIq870Hgrayff1GnGd
rQgdFKtuWuVEbr045hUZBxhKTj9VYgOoEyhKOZQHh/FiLMQmhzo5WaMBZua3PUcrGQYfz+FiTii8
Z799CNWhrzguE1285oqMLy2/82mT1NF/HU/WbH5cpH+8an38IuH6mjp2WQZWvBc2kUI63cU2LMD5
8mN6xpMftETFgSF4Utw4DNfHFcpK752OrciBcqo0V/TOzirrVXmZXM+wdboJwblXKcn4p4G2hgWm
EzahPxaTpsN23iXCpbn06jJU0dyN0TawqNutsSg+bw25kr29hv8m4kr+3gnI5NwVCuR16vx4bdVM
qJdJu/6MFgk4Qd1bwqyj4UKMCt1Ko/mCeDA0ilFS95M0kVW0OugpUYaF+hmOIwmAOSu/EFEzP62I
iA/tKRopK6bWu9LhyRM7IJYaRJlHcYs4LtXClgArtW+dx/EB5Jv2w+g2HI1/cV2wvLUPDikp7X2F
g7qAE3qVcCtzRih3b4qrSUNkHjPFKnPGbphEXerOmxkVxM/pCfZzcrYzNQl7Tzt3Bbn4JT8LXQlY
7NXL0r4UBS/Vr4cPC+A1Oyv8GAeRpCI/eSaWd8PUdBKjLz7jAWb8/eW3FpWHc0hLeFqM0u03RQBJ
YVgkauDJKVDHfE7K2ih9UKx5+MLv5OlEf9gZwXw77flZMhhxWrr0yumcbXRRPHhiwqPmLNoK89uH
6ZBixxQtbmewsJoOYd7QwvrW8OffgfTOhzFVefZKJ1dRrQcUkKXdnw2TX8UK6Btg7TTS3vTA6s3G
lbb0bDQUlxQTxjMF4YTHrbvdYqDWAYd7nVbujf9ejVh/QrFGezhGZyi6AUK3U4xNIyORWBeu/HgP
Eq90sR95aFESqVZdaUxneapuRX3+IQa576vul66mHehmtS3CeiKg2aYyHoiH0uDNeDmgAZjacmKc
stpneFlpCj6NUWtJOj0Wntl8oJvIPqF/1L6xwH6sGjCCiXrRfjXhlIPJfUnSIiN60l8MiPjdRFjy
rzGvWIch+zntiYL3GzoxqHYriCAy+3cJHu/9tODcIH6fDJlYVsk6aquW8ZGGUnQ6DDNTdj86X/Wb
nctFffusn1GhR9cdylccKSvIxhKMVNLzIr4nq1/Ahp70vEd+TcroVamt5ofdUiYSJLAbueSB5Tn9
ec5vkbKmyE2oF+BJd9LTzPzVcScV8aYoMC5jVmiO/jkfrtC5Du/qVdXWbGSElDAgzb25t8Xt0GfV
5CQDJdH9i2mqM7u59t+ALkCfvLPYL7XBguiFD5PH7o+M/9Et4WbFjEFT+AYdJIYD61tGvqnd02WG
DUHg00mu/xyr3hVrZXfoZEQX62eQ1NfN8JcukkStl2vfLVGlgMG7KjfbRp+7XfrIUQvL1qdjoAOB
u+PA+jY8G4iBblkkpbvYIbI1CtjxuQgIMsj3UwpoSfaTtXOPnd6nbXbRyS7TITaEcROKFotzpPcJ
VO0eoXx2yq3hS88Ty7xpW20+1FT6Good9bG8u3ZBDf4khIbsybBvo39FIRiKF+GQRSZDtNLLrtpV
rIl7N2BwAKuo2tiP7goUGeaA41FW/i5syxV8xHXrTnaMDtV+27MazJ+OxsfK6KbsOJ14FqFJz4Bi
KwuOGmv/8V/IBDu3+rpQnCkcc5qptmRJs7rm8Lpnb5FInlaZchwkaBeVnqk5CZcGJ1bTNurYyyvH
xdA6WFafgrxpYjXBbePCuVaH/vxNTbHvWif3mCGKd9owvkSOt+RGI9WW7cmEE6XkZFevxMid/wkE
T5aFRh5SnMU6OG05AxbK6IGXrq362DAVwYBRwIJDcIpj6/UWESVsy9k2bZHVjRzy8uOy2FzBW2Xy
2iMJe4H4XPsx9K4oVnDUquojLttKZAez/S2n5VScu9vqs5zCxe2QoHXlklZ0mAKh4JqV3GyBU0Qv
5pHwU2liASy7I4vvvsn/GV3JjVvDrqFiiBHwofFYAgWSL87Vk5pUFcBgMmFa/HHFmNBjqq86qj/7
8ZKRE44mhk6SiDNKTeddKFTa+PyR7GGscKAH2UaJdthXs1i4B7IknL6VIdZQJ9nEazLZjsnWhYwY
RF7VKm8NNEIDeUyRGZE5uns5E+5oPhWY7/fFA9WER82o393PthiGpgE1lEMNGg+Jsur38+0hgDXK
/zPr7qbfmtQ3DsxOfwObig9ha7BZMiT7jzwGl3ovlY/mGCKUGpnZlyZLN22Fmc/71LMazePZfu14
gpDoCWamDxb+whvmF0igAsFWInaIiHGeD9M3ybQ6c9ResU4BO9UWIUmAxRoGIJFYVBGQCy8SEJdc
Fs/vbc9rYo2P71bhFq2JEwpJGBEhuw1or82/sybwLB0hi3mnwJNB2OjEF7U3tH49gSHlahGrqtC/
X1BmJ2Xc1UgHdF6PEDFORZVfuCaVCSYt0i7rsvgZ8D7g2rzh+AW3tkTyppAnnuyzB3JVz+lXP0VF
R9HyCYZH3JZWBjDs1+wwVpwCEr4ceLYm2ojapf7GCbT23L5imNWSQ57XDfUFOyRIfdjSCNB7zpuu
WgNC/2Sv7B4FGHDiFcnGuA9ZAdKxaWIejNPKQDRXZGXAGSMDj1GxwB89XHHqOCDEf12CaYIVTJh2
l8pZhk9gFSlXw8n5e4FcH2kDJ5rk9bNblnZFkueHkO3roQ8uyVdy0oRXWJeVMvZPhoF+lQZGl5tf
ADryohn0SMOYbBLSCm+4Rx+8YOrAjhTvDBO6C+QQ7PxIUNEsn3wLSAslbvPF8/pePhqbjB8jUMww
4bK5hzVZEpAl1qCz68vf8DLS6MvDxB6pJdmhfdMiUZB3EiphJ5y+RF4CGLGZj5G0jvld9UTpMJIF
tBfN9rBL1WweBdgmxWD8PQgfUMFkNmAWwOa/wBtxWSj6IdSZboFoNkL0iPUsxV9ufphVv09iU0PT
xQnIC9KAabqRuw5CLvdc1X/aWVPZbLtjYVzWnwLE0atQ0gSnc8P/waFx11p4nzYLVt92xQwLL1jg
Xx9CiqWRLUo+b5KsVnDEHnFBM/vGvP08Yfyvay/s7620hqjJMVsaUAS9lNLwQyHh3JHpDPie3rZm
JdMmY8f6UM9ESLjjVooLVb1JxXo/e1CgnDEoPdUAxSa0hvkFF8MeuygXGnG7/i8rRlMk3/6CQLYR
MFTRKoMlM9oS5TyegtuCw6abb1UenWgMNST0w92jqHNSDmPytPUr3YakdOjIcZdaUjevpiPEMrMr
cWsWHWowglHYSf6pFxPKdi/BMqFuJBKCCYJ5edllKlBb9O+PKYbFYE66XIWYYks3t2QZ0HoVSQB4
p4vu8l1IkjxXGKdZcKK2FQkrkGsDAXGUWnGT5E4J2p3t4bTmUb47u8nTif9qf1ME9mZ/FLbjUH22
9g7K/MDnOXqE5CcWKI3tCzs4kT20XnLhNdoTN9JEBhtnGOjtcCsK4IKOiDCtbt9KvqVhkNP1G07z
VOPvM9jTqFQ+OcC5M1p4sRLOT2b8Gd6oLkxnHt3XXnPUj08uqJkos3BoaQQ6MXI8yOREnwmr35uC
xHi7zF/DcLNpc1eD1n3/Pi7UNElKxltqIVYGr9kwfQtHmrTZ8qkIWBxYJnU9s1eQKEir/YdV0/Hb
L74V+n8xaWv/vFSDlh0C/hntlUFKWhVIcOrfT2UmCEPPc84UJb9i/ktgv5uSr+pxvAEt0Lg/Kg94
5VoMt/YzsmV6Ksv1AGIgKYGI/b5EGMQE2n9ZgVN0W/mVT51xcGl/+v3WlPaYFBCBI5vX3/LpRqon
7c1EqaHtaplGduQ8li3c8827Wu/MtoFzUJqdU+hUHt5SdiTVLWbRCdeGeMytcKBD6ez+01FZhANt
Gj6V2eJfqgheyeZIb9wrR21D8aq8ZpyJtjGPCQp3BqRNeVAAVhwaCZCCfKbX3oCxa3CcThtiN5A+
LMtFlun69kSkbbpQHRxu/rdFmQ8NrsquOPyHMl/12dmlbTIgpj1uQKJIj+dJdE2rTBJCSgqAINDc
9dF6Z01IcYsZLcNAKzsfYHwuNp1KI/R7ddqBi54vMhGC3/IlkrPVt8v3fAd66NOGscl6jKKfPNFK
yqUxT1C4i/lrKlZ7yzezRHB8ZLaB9X7jfQbSopD8jixMFwDOmZyiffJtTevnIEj93DeC5CbuZREP
EKRPLsPcqKAe8Yn4diQ/01Y2X0hTy5tE8qP14EHiIQl1BLB9KROnrN4jpPTnenTe+VA3WNHTY/sy
MNQaAnSkh+D4gkn7TbI7mnbqvjUr2t0pAkBGy/eHsPy9h2Bw6W6qIwhZWyWcOSd4k/QaJjW6DiwH
DVxv6e5bTloX+UWEUWuH9P9xzWONs/qUEGROLEClJi2/dPsZUOq2BHDlcfTIWydwrAJBmEWxe14Q
xwFeNkffFkRkZugu2OBX4RAYKup9OF5yzxl2jVGxuSYknckuJveuHZLiQTTvRUhRdGQp7g2xbLVV
VfdMpt1fpKdLggPyDIPs13FVkhKMXq+6fSE/j55DUoA8UJwFKpvlq7w6kf/e+lX1BJTGjtbTl8M0
0FE6AA4hePTY9ZJw3ZaC03drGIl8ha/bj7lZvA9m3gAOR08VN5gfGYPRCIjVpTEmFP/UJlF9Lk7x
bh+2G8zceQ9dfBXuElfbG9z7cfDre2MkiOx8JfdNg0COhtjkNLxDuyrhaVZpz583LXYt4r0wCR+R
9DEU0xLjx1exRFNtCkPAZdKzA5vWJ5GHjOxk0MlkGf2bc1CpgTSD6CEcUrlErNW3TxFYiUGROmAg
hSO3I58jHavAMG4kHBFd0EPtbO4XNGURcbCAlMUk6zoqQDRStaIl4BR7OBdJEll5EQpqNulvP2PM
4DD4GwbkFd1Npz2l4LC0sw8a4q7nfXCbSpfe9j3cddIfPitj4kBaAuWFOiAL6WbVnDhaVmK7wVCk
AfoA+YjgWrFRxgcWD8lgpAiz+Z8b1MAefWAKOdjyRUSNquLlGSnu8Gdhvd14N0fcX5pryxkPTDG0
I4DnVST9ATNYdzEZlVAkmEX9HSs8c/YYKZwctj2hK8p33D4u/vWPPtA47QZM6EoyZahtb79Hf27E
6e5LAY+b72yt/90Q+5VCrD3H3i+zS2Rxlz+sSO6jJioYPlNKx1BWyq1SiDaYUVDbXJBgc2vV3vJV
B1F/ao/AJM5f3I5NpKsZouW6mNHY2V+uGTtvn3dePZF5OZ/dXwnIEmJ2UQH9UiawWXTl89fEUB0T
4EC6KfOPs20xXc9yfjwqPtXq9vC3b961yuQmzhJ+cBpBtmcLHcd9GGtkdJ+mAisbYANtBMIweavY
hswGUuyQNbVBcNB8obzOC7J8326oNo6j97DCJsKjXvdglfUefVYUVWURFO+EDAkv1Dn8+ciTv8Bb
rSDDCN6gVR5hyq7KWKdAS/9a6bZbjxf/hLMpfd1KPo9lNfIIdecuPnXTy3n/3Vk/XkrckG3tqB+u
rJ23aPX0CyML6iV9Ct5dF0tetQxPpMwF0ri7SjLfloHxpKhbcCK9pUenbz/fFxagnUIPWXyU/YE1
JaB7yRoJaM6TEn9rnO0VS0FRPF84g4ndeDFXeEsU8kREI7dkLP8ds2HXzicT+d7gFKGDJDnNpqOK
tpbXRtc82WvsYweIdw5ndIAzFExeP4UlOnjqiBGdxAqQtwhvjtzzKUZceaMEGKxM+kq0Jo8BseXf
8+BgMzKbfdtNCFzN3w2ONqEazj6cixP9PvMnSfB/V4z/b1qXbBPhFNKG3IvVM8ZgFdmdFNBLivVJ
zDTQ6J+KbqVWtBILoHdq7n3vz21I/RVAF6z48Zoxm6YbW8k5yEpiMQgVOcQQQ5FxQzZjspvlwb0K
TMxHBO+xm6hKs8pV8WxIjStM1/GR6bIrrBEEkK4Dlu7en6Cczghouo5pNN4gr795altOU7ceERti
mB9W5MF0pGYOLaOf1LMjp8W+qtb7WapSyORj7ahg71qAhnZt6I+x3Son7OAVzXpJYTrBE2nwgYOx
klUbhCo3tGnO6+Pd++KBh8/Wrb++Vix/quBEm/FvTdWxchbxyeVfDumy+8NL8mem6L4npBR3MyB8
3Wp994imD5VotK7d1VhmgO80LvhZr5kTPiFl0daQLsJpbFEXkz8VDklqIFSc0MHL2MPcKDhdWHcZ
9XJddim9xvWAcssdPoJAog23loVqMbF4ZtWk1vcGn/Br3KU/K31TZOjlsnnGwpKbWqn+UQcRGmaK
4yUWdDsN7I2SwQdNQ3bv9x4Sxdwt+lDsYoeHLUc4rWYfNNKz5rDCMQvYjDmbTQQcYR6S11dRm5GB
cMVAm4ngtgYW833yKUi+LVyaqzBGRx/2IBoKIMtLINfQYB+lOeMtBhP8vK0tFHsIEwIrWcL4kUwF
wzyyZkNR8m+Qs3HxBTep+dda1PMjEqDlJRTE7viZyFqOnBDvD8SRMGlEDtHnzv+MGx6WiJ2FfTOA
vFkfIyg6XX0O8KnUNz4vyjsz4te47ytcjzwMa7DYlc6IduEja/VLxNZqB87v2HpasJQXFx5ToSyQ
w8yRicn5/HGg2cTBTHQpo5iUoxCBxDN7PmCnOO7zDYzZZpf0KY2deuBDNt5TmJwJQ83L8HZ/sKlO
hRNgMB4qaVfcptgzxkDqtn6FvKR7IoJmIGOcWhbY9wjXWgAkbmcqLxhZAs0YQV1sVhouWHb5Qg46
nKIw70xS9puPnEJH/kKOTehh7jABF8x8SCk80WwggG1BWGAH8+D1CsppzLcX/lslhvUZN7T1H4a/
LUqh5yvRHFiwzBquy0RQcgO/X2vVUq9uY1Dkkf0NTQ8m6HKOM+7tFPtoqeKt5N8Lvg4DRjeJB7bg
V6en3StC+tueyiZODVioSyt7lGET0IYHmRYYMfQRezAsQPBfEVOga6hLGUoUD0r0J0EphrBjLSBq
y/dR/osrxRM8+LPz/OabIYJdBCde/phL2GmIwbIuq4l8HNZyvn76nP+GMjj0IgDt3Q/+6jOr/+sI
tgr13R+B/jT+X15npuPYruCzW1CTIWRIEDPncW+uZq14qvWv8PWwPGPtVvM/kvS0wTsNCBhm8O+c
LS1Uhe6zVtLt5mYAVF7ztEPZ5wvHWlb8++XczT6zYBdvkGcbaQ/YRaJWrtzt/f4ByD9wBA2NiJOg
4MGR2hgjjtzK3NWLs2lSziGfj7FXv6yyLqo/Ma0yTu77+BdwNCPoqGHZQoKgbiDB/p2EsDMj9UcW
81qYuCLDPKqEe0TrQUXVWvfYFbw+dCFMqXYAXYDqYPRh5rSAQior10rOazxnRifkDUbXiPHP5qFL
aGyDmgQZJhBGSLboCu2NVTKVHHKJ6Xi8IJHGo2EQmZwE/k/sNVtibKbFqXVFGO4dB4dm5lDPpFdr
xug5N1xAHmrIELfNCbVwMM42IJNjNbPNhFgZVAjz2qO4sPJuRPt6uqRRvuNqkxWpch6b0RuurufU
h6/Sac7IoE0O/XcSvChoPjSDe90EDwmHsUjdZLxysLVxTuXqKwr83Mq+subHz6r6uf3sLJkjzPLX
hmQPzUZYcmhqcqnCDH0uc44DoZ/Eb9fA0262EXflOYYX59OjBjoqvkmluHG9WUI5waGc9fymlbpQ
nqMU8JiZrgEkjT8t4FtFwBAWyjPuGjOj1LT0GtWzQDUGsswr57eKxuE6HRIHHc9QlOIXLd/JEwx4
yD1w5D0gfvhbge1/joClQ8+AO7pwraiV/5dmisrrfty6prNLJ/el+ubbLuppItbZk6Md3c9gOVn8
m45XuDuh7X2c4RS9MZV4JHVsUo4gZemZwG5Kr+oK7hK67hx+HaSXXlUkqA507n4z/BGGkQmnBAVc
DZj122lxo99NQH/N01dPhhUW0VaizaCwq82iyYZlIjujSnLlMGi6v9rTydyRi7clAN/VI0ouCS75
0NaS3LpREqclG1GIzfPe7W4CNHim+px0PqmSeTLjPRUMDuN9USe2sos2cIMNrTBcDup4g7j/RPoa
xfoagJ+0JpN0dLnqZVSxo09BQplvZaI8RRhZyLLqAoEO6NmcoN9WBObsTSE98Sh+kod9p542Rdnw
ueNUIHFPRA5ncGwYJ7Ko9l56ibSbX/XEy54Cu4Ekm3MALP3Da+2wFe24A7o7SzhQAn0vfarhEg1f
3pke2vDPWsx6+H3x3hYy9B7eAvBmTrNI4V9s0gWBUdi9JNgnHMSw/6Nz980fTDN6sciNtnEo92nB
8e6Iz23UlQ3d6kVbmfdGzQAJcs+Ke+1TJsL4D+x1IxqI8O01rXV8z0hTK3K3pQr4MMSMl0QjeRdg
pwPd3E2neoQ/aY0zksBAleIysPQoIgIl8coAONAw1S3oGJTAY6zhsqkrB2gtQHPsg3aznC43OyKb
z77e9s+eBEkY/+VgNRHg1AooYWDSLdzm6rOuLyWhw870NmBswEd+yvjyXFDyJE15/0hoD16DUKrh
6Y4l/OOom3fhJVDrbter9TMBh53/UAVsH9OPuJ+3xdoYa8jc0POuUDlCqcDL9+rksH4ydF/oNzB9
K995/8Ezi+F0toaJpXON7OR77j/u8diSeRtrS6N3cFtE/zaQbw1HBOXVcsyFbsIYQdbQZuuLkn+0
Q/mrR1hyx9Rq+y/gd5v9iXH0BpmnSdbTpiwJHUfp8LNCDMcXj8xSGWqtoiQTLIlJoD37WvwOv8Sw
vg4AWQc75A+zdEecq1pzXm9OzE/PzRQXPz5qEd+viBAVU0O3I05hRYv/yRUhukjLBygBM/JMlTTg
7xaZOA7ov8jl/BQ1SqocS36i423/WP8m2902+zLLJyq+XyP2OoAurLV+49WdsYssimdaTR5SAXWy
TF+Hmd50W74lhMZNsglJE9cTJ2SCT9ciHz6kPtyhWKdLUknjfz33dyA/a7wJWTDUF1/Nc8T6AJhU
mocyGkkk2VliZ3MBUuq4TsMBxFlLOoMNrvLTcCQBywrmjz4WrrBIf3KWHhmtsitH7HKO/SFSQ9fc
p3BoRkdRT+xWD/6zLSTTsRF0Ua/x3Ue735cLKtdkWRDQv75fNJfkVRRv4rNIX82QFJaJOxfhRnvW
mBfZ5ioKAy2vucYrEg5ay8S84xQUz7asP69pfqhFQPWyrNZO+pIBZ5GbPyiw1InBPKdHfVE29esS
PcK+u/t8RfqjixqbUQGzJ0rMHK6XWeUEb2adpkousIfXriOrFZwILto+ZzbinKNzbnlhcy3re1U3
dKXVzWRfxV8mG6MIduLMwrIVT5MYzsIfAPnuRYiGfcTszQZnuoILdExzmrS6S9NJ/3uoIMS7gaD+
Ih0gxMYteFsxXDrg1g3fJzwNkQoEBSl+3SsQt614qFOsrqiBcHDd39PVMlQU/VVwU03mtZdCmS/s
vXdpuyYwKFVq0J9y6wSTZ1TTAoKxzFRO4PSs2Mware7cTjHRUDp4JD1M2y+kJlO88O6WaAQU4vrt
qDl6c+PkFRRJN/EmRQZGxi4pQ1hUsoY07gNo/iunwwSN5jdAS1Hu6Sa/DIFZrlayZR7IfNHn4d/Q
XHw70t5O1lV+67WRI3xvWFYs+0pxkj54aw61wFnLtCpW1CdHPKchIJ1IKgfCLQRu6JlgoYI03rmO
HSMrcXBbQT9LZDg8sTTq2EUFSWDmsu+PzfzwxT10Kni7eKOn7J3kjOH7yAQfBdCL4TN/5u5oDQ+U
ytquEHDySlrWUQ33R3Zqkqys1xdtxQLyMkgjj2nYnkyUc/QgQzf+bFFMFvaj2n9IncS5TviwmZae
U0LUgopIh3BW5qnv1kcxOBuqvNwU8ykTBKvA601aOrrg9Ya4J2Xm6nmwfwlFT34Vrpop05fIFvRr
j21bVY+nZvnOQKW7TAYVY68FoVP0XVbhN2dK1H/K1aYJpntRAuBLMpVxdIYrILH8iIb01DhJboHn
ASJyPGMUYJSvKIk8RPWujffQ7TNVp8PBc6UhjbmpeeZpCJmE3/UqN2aEsi5edh6DKBpbzj1Rc7d2
p6oED1YpK0tf1YFwjr/7NxIwMVKwxDX9quwZ0j2XwHhCRB8bTghIs+qkY9JgQVU2Ew04Bt8AI9vw
i9tEiJiWT3qShiRclsbokCUAbulVv/Dpi+BBAh6Bmgm4BTJlFYu49Bzg+C09Vk2HoIKWEX/00Cas
uQIJL/Vtvm7m6cuj3hfWFOzc1wZt3DIyYPdqVe5bIV2Yge6B9QhgRTqbclv89YmZDVmknDsvBCpc
ipf83bpnvep+IuTK/ytvolJBiSfKP7ehyPyD2T/bt3IZ4halhIVmqqUkFHHHtXWeVm/WkXHUX9dK
02g0NnU1bLRVBW0WT2XyFubWGdlKQ+aUEDX8fNp/kLAARRpBOsqoImeWCxObsy48zpB7e/91KQtC
FnFkCTcN+YynwRCncyDSLp4tffYRVaU02k5T83z+3NArMEwhe7dY34d+yrT2N/AgNohY2XTPqZoN
UkVGH9DWqNiI9DE4DrMUs46IyTZ7rqLXnsSokdd8m+BFEqI+6h0AU40Lh1ahVbiXjxPRyk0ZqGSs
km8m/vi6zCmZKJ6qq6sNZQ3SYlXQ+yk8SQN1pc+gbpm9CLf3m0seVewC9s28yqImAhIbyP2h8bcF
DuB5jLPBZN/NWDwPhaUnOBtj9GZC/tqmVZj+v7Quq8Sd/zYWDMMU/2ZlJsW5T36Sd3QtYjtlTjSm
+EYxcnkv3rp5au7bU6vFSNkdtOJ62RAkAysaFll3rxQkW3ehDezDCBNYZauxmwtWAntq8827EaQB
9E0HnEwKQlCzyQ7WhKOVss1nu6ySaoEGb8wyIusYmGkGokGcpcYQ5acnZ+MIeLB8WqJiZPJNUWCd
uFYnWox+z18veskua1aayE/eOAZku7oHIsbpTZRGAzetQXp8Q40R6YwqFrH8fPCDrd7TERqZ/zyJ
/MFoqH0ITa9htYpQxoJJhYEZKsV56NSQJZ68FJAOd2T8Gn2LGJXkINLJSHbk2L2XwKOhf/LCbGuv
uN/xsfFFxx1nqGifhFcNYe9NHrrYmI3ZX/8OgNNkLy9Ripiub6Wzw9Hm2u3Mm/LkpjZDQQWtMuds
vV3LX+LUIM90Djh/zNmnzEkO6doXjLIXJhkIFWWohYUyyEt/rWUTB2CKOgaxSCpObekmj9zmOYAV
eniJp6lrbIStuoupIdwdmM0Me1xR9cq2cD6lpq4eUS5/BZ3NZ6L5DettVg88H/j94CelZSTKFzqG
tJVgqwVk3S3X3vxuufqTj6bvqdWs+LMN9DBt0gqL2C0myCiNau16JVJ8SBirlL6kzBK7686vPBTC
rmgmpU/bnyNnzzVrf1x1T4/FPlcgdP9GHhanA+OWaWiQ9G4Gb60BVAsOtD5J62WJo+eWtkrV50X7
O6ttjBgk0UZgVxH+X5pxrg17sBX70f6ufb7rnwKiO04elTCLncAF1qMny7iQ3WbED5DAqmiY2GPN
SXCd3ywSCQJgFz+QfLPxJ56inOpHnOQoh5k5/ePtrFsAV9j16JlYfiPZvmmEDUE3/tj0b1gR4ymQ
PS6k6JRuYkktJ/OzuxeAdsBE4WArXyJbP65RrierBfX4BMOy5xwNJL/3lmG5CkCM2v5SxIVe0RIr
7GeunSrD7pxEq39tKdMj3ttWxcxM0A4cIv9BB+bndzczAQjuYBNl28v5m6NHO36vyXjqZ7aXT99u
3ArXItzY2OpnJzNf6QUzSXtLEyvNjna9v7ZpxotEXydZm7P5PGGSAJKVSZsQg64ccGbVzToIpX0D
i+0/yJ+xr+XHdbwNDOFSjfpYndpflEZjixeM8qbgzLgPe+iaz6X8QgBF3CZIgOvqgjIRm1Xw5cr7
8Z+7fBjQ6Tz+4q5Xtb06Zu+5/rGzNojPRBIBIqL8nJqHPPdR227EPNnmrYdWICTuvfRkVFPEdnnX
8DcreMDjH44Oaxi7OIVxMc0u3ZnBLqQErFfsVNxGGNAVsHpCaKrrmnStYU5PDHp/KdgZiG6IQuIW
gm2qfIL1lM5WyrSs51j26/DX6g2ua3YYKzy7N+ZvyQrS40koYFKbDTgxMTqUHxhSBk3m8yTZnK7Q
Fxul+tGLTfE0oElsk4O8gG4Kr72XnRRJL29FVJil36o6SrGFtAkqXwmrUJ4crwg8hcEsNtOaSkRD
GGB/uJ/brWCk4v/DW5u8Em2McEwo5cSXKUXwKF5o/8+0snebe/O3Wm+QX8GqImdmv1VcoFUwoYc3
SkhGQK47cNWiuQRw36JZtqg7dZr/uq2ZR0WpFQRCufalY0UnmYqWetCh8MYP9hkioCWUJM8P08Qm
nDU4UmC/HRL97QoICaWP02hiA9r8SspDltYN2BR1cW3gcaVdQfV9+cxNDiFvKLAIZqKo0TfKCvlA
4cTu4R3ndUdeizSIFSlRmdjGpyHC0A9YnCh6IujftrL1ELv3tzQPee0TsdN3jlMPUwhwaQXA83Ja
vfHKP/eFZOq6usIFP195/u3O1a6JbdClXa4AAb68Y5RSgvRHp3vM8sQ2gOMVBtKDEPy9Eq+tp3wO
ZJWwXhSgxTdDbp+t2uDkKzUgOR69bKAx9Aemi8xgLLauGBfJH9Gsd73f1aD9TCJmvbUrSo5tOvpO
iD6iT1FyznYqJdjP8aOWpLkiXIVrn45NoEk1pqOpe8nz79govnWsIJc9eQP2LVmfFBLvcXT7VQ7n
oCHGhehhLRo3px4AxgAguGY1pqYyT5krD7ns85yM9ksjs/jWj3rb5TeAzbAp9hsOAChzWqlTH22n
DLaiMgQmR0tpECpHIJWWPCizjoA1M/sH+DEVEeq2m2S9fVwwBt1RifEibVSoM5vLFHu8EFa0Prxr
d2EwDaPLqDETbCVtLMjDHuoxLQekjxaQPn3sDj4Op1asDiLTyvJtRpYCiQ+FTLX5vnyunHxT2F4J
uLsMQuXwu6Mp/f9eHEYQfzIxZuMdaDiRiByem2ii6npnS+/00us2qJJMgFF66B79BcSU/cTH28QU
wBjP7dhmzwWwg/fF5DJlT6NWnkfuuN34JD9OxzmWB8ZvqFah+iVwWCAhnE/j76asDqiO+qBKsCMI
dHVjpHjoSXISMEinxt3GfGQoWyX8ZcXmgoDFsl2yweCNfcNjkc5YooF0UJXGQeYS/emALkXsrCB6
N6kIzq0EGIjyO2SJtbLPSloTqDs9fYDuheAPB6rFkp4+cAsZyscRBr9bDu/rxqtsRO8suQKB/IKs
v5RTtqBoDqelW98lzG1H/U81f1Vd7AWjH/ScLVb4Z+iMRod7njA/KN9tLSbOjBHyPGV6AD82vj/p
8IHiKZ1T9REpNGATx24zbe78P4uEju2BPDl+BPsFKYRnu/9JPsaXLycp5CPavqzSOmX4EdJPKLnh
sncyJX0h5abcCzZEXOdmx8kBvsjXyk2F+WhKED4Blfqm9mKyBKULDag+K7XIUBwg/54c8UEcneAh
amM1N1WDjkMjlUk0kPUQuvjzb9FZf+rrbn9SqHDreMJrR2YIms9NMG7bPopVAi9MmzAIB6cbDvpN
I2SUJ4VJM6Y6FpScZxRsOr0UD0RB6Tv+bCnu+BrzzTWcDSkR1sVmuPUzIwd9Nd6vmnCsptTz1H2q
fj+KzghY4BfM9333VlrhNSM+x3wzkQA5+OhDCMKLD2njoJ9NdvQL7UGpsNYcCOkX60tJNx0H9crJ
4Ze/V5lUL3bwgEw/wEK0DO3AJVepJnkFz7AewY018BT++pO6QcMV5GR4L6UpVUAfVi+Hl7kXrqcq
77GHPCZVThnUBRxuwE0I0hAqtl8VIZBbkJaM0sfpZ5qG+v02zRmgbQ6/MWZP/OphTZy8ZhOfJ5QQ
6Xyk4OzP2WLcYasKUtc9mtJb4PHK/96s5kXd/jmYX4Om70TNCNL8Z+SM7L9Oag7dS7tLHQCfqzfn
ZOzKnzdkoOftu2hIzFxkvMPtP0R0cePHV4bvD/UvoOLnNRnaHYYtg1zozZZZkufHDCJDG5u3OBxh
imoDLzRm2gb8kNRNAcaEWQK6SLmhxw7QAzcyg5Yn3ZJSTgXkWYKEK2PuMnlHxv94geMZiB2MKV1t
jD1BGOIjBx0UOl3k0ouXkQwmn7ZpkflcFUxpf63dNQN/QoXI6F+ces4Fnk7aFoVQGKOpW1dJY2tr
09EKpvs8Acsw18+s5FoAnjZvhVzw0I9nl+fTbI9Xx7CoyWEhlD3HELGZ2GP6fbARe6eE+7asUrJX
yA/tbb21F3WjP0g27ddw4LdGDjmA4dBWEJRpxfxeEL8xqvgtTAcx5Ka6/XvilfyPkRgZLsYHBGjZ
NRTx6rS4DCl5TYvqQUVxYtRQX7Sd0Jfydig4bPSqW/HXqTziuOJejoEPiRn5ZrEUdUCGR5l0DAc+
Y40ajsxhmaWPpnJDKdVoR/6C5U07WFeh2Bs/dn9nRwGyiXobP4oQLuS8H6adrG4vsfCsNcKP5kXX
JwxCyV4RrtNvJeJoanpeGKcG631vrF4zJ8e/+hFuvgaYPxtP5Ulmg7K0Sr9NC+oX1LLsTuJ0buTl
LqpSCkAk6UlALnFpiO111Uzh5+5hkqr6QIPpK6hsfiak325uC96tga13VUOy9q5qGB0JiILeS07O
N2tRvRTk2/rXj+UfdYNXLhWVh2PYPJHOwBs2iRczIsc4OcXxCaD8DfFJRcIlFa+W6gQl/SjuyTKK
FG2GXsgaf5C4MYCwayvV5TBUCqZklXyu3sgWjY2WKdFVVcGka7+taUQe7Z9qa/xJVhGFe39cM8jG
Ogj8xQbs21T/tFPy1THKtKSXGQPv42z5jUs1QE98rqEEsK6xW2WQcT/ZNELw8AiIcY79pinCt3Yx
EBubNRf/mM9ChvyvdJqn2c/IC6fNS+7UZC8YmG310qLF4r9EUVFDxB6rZaTooS689YS1IDevkqtk
ul7k8JEe6e1GuRXRmeFVgnRIXV7bOV0mPQz3wtA/YOcRKHSrPFcZucoZ5zSH/yD0U1R5i02t2TPw
CQ8yUt9TyVALDTEZTg9NOFnmzKxvceJXqcCgmhG65WKGRGGmQCWhqQyKCskIJ73bQDSH+dNWpXxW
YoCPOYqtIzSRo1UFFmt1pHJYUZa9/fPIEd7BaAfCCTzOs3LwrEjNEcItaTLUPPpp6cOwRWAbk1Vs
2Hnt8jn6HKFpJ9UsnAVCEyQp1kXvkgLDUA4icIEAONuid6YOWVYnAfTnhw32WJ/wuwaPlCCQMvsH
9dUgRnzO/M18kST9WdxTABCoxZFYqCiVkMfqmLpm8WocXJk6rl7vAN8qbpA32DepWQfu0GOTueNy
9BYHiJLWiP13NVLxA6Zi/8vfzUUbrAejCiURdGgFwi5F/1su27vJl5WgVzaOfJG2gd+7zrOJdVCF
XZ5UkUn0tcDJW91d6uYShOMxYAPpO69sOQFm+/0UPalg+ZFtaQVcCv3h3Dhz8RQc1QOCg33zKB6z
NRTYiBvKlfaqJ7b2HYFaWr74zk8/xaPkxiPFdsoPTCL3Z3q64ctuSyARm9/R/gXgUowSBzgiD6IO
VHcZdytY0kJBuDZCmAGUuqEcRWmjwvmhoIHBw7p0AQdFtjsSU9wSOT08SJjoDp7dUhL3eONpC5w6
S0iRWIsX6uv4mJ/jcyM40T/gmMjE4jLqCQlTz95BGxegmFs3pB8uQZtL9heXfPbO0m/PQrgPXZ74
jNKhBrK2ekE0pFB5NwW1VzmG0aaszwAA7aLUP1U1iPCRGjd79LW7biZhsofzLB2UPwwlrp656lwT
Ovdc/L+HkexJtV9KNufd6GnDhUoyggyydqN/9ALOL7tYkjviZh8htc8T5iiC0m/e1ng5LPC33GN4
yP6uFZBAIeSi6/9wA3fFsF0ZDcPkCRe8zEOVv2JnTXn+guwbQ6sAhoMRDUv5s8Pb9mZla8Jm3C3G
CtGN+/FaECvZ7d/kqeooIYBW8os0/aElOA0k7U9p9RpaV4d1DQI4RTAFjhu5FaXlXAsg6cPcSRC7
ArVczLEd7vZsflJ2IcbR9J+oVtPshVQQ5FVkHhQecCNmW7MXiDOLcxBbpEvQvd37ezgiUbeunqEO
d8Zs3Vnq13yH48eZlymjwd5+Hbu5FbFchoWq6Gtb78Wib/2Yfw0YMo3kmOP4sqheX819085iX4Dz
8O5G9xyhCOnkl2gnvcDoaBACuimyoigiTqfaideoIeez8EI2mweccLR7E5fc8+GdFFb2njL4lczo
IEWZG8AIsp8yIQ0+i89pwvKetPy2AxpX4tvgSn1Yf3lhul0i9Bv2lk03vnj3amd11YxbBAxTJ3/y
ArTa4YVR1zavtg7B7crwJ/3tS3jI7WU21w9OY5sm444P5hCJqupjAYLS8JtDbQXUL4BRVlANpMus
SuZEY60Qo35dzmTGad7/E4ANuGp1ntoF5ITsc0rcTu7Q9o7KdWALrVvyPk5udF55yexuZZo8b5Id
9NviWGLCiWd1t7zgsjSi/xa1rIRI/ViaxzPuxg9OzFWEyyqcyxWHtLxCzIvGsaoh0toG5dq5sVhv
4ZPTAQbAMk736IzAM36iawUSfennDi9es7twts6zIKzSKGLBvcWdhhS/gWGr0v91mVjQR8ywxtD3
a0+7TTcr9Y9w891eGqSLrymBjXRBTqSxqVt8+11Cy4TFxi9ArUSWfA5DF2coTq9a/xocWiIR+7vq
tJ1vhgm6LZNB63XZ1l0tPQWQ1KVKPQ4iGQAdF2iaT9xVDu7RTL9N8s0wTL8a2jniX7u4JEvVLAE7
Fr4RE/RVaeaATWgdkgyHva+CK4w1ru0jLKMXFacfhWD0OBZMHtHmIQDsbmPlrTU4vWwo/LNDNpy3
s3ognA6Gi3fP7tH7yAyW/AJd6RYvi3o+KjQkLF/lwNu7dqiomxGLNw107HE3hDA61Q5lUsKfBqRi
GsQc48jsotmoOAc27AcdnK2jmwG5mNYAi7eoHpHpJYIcEkCQyNuG9HtgcFJoC0OYkl7Vn+ZKXl2g
X3zyAwBJkTsjXX/MNMtM+YoqGcalXp/0WPGZwsqY2l+n5N6pAw1JihgVWzvwaXdSiPL1qgcV+MQc
MVOP7am2s5s5EAuzbk6tBiqgfWBmMEtS8myRJYTXcBPTVyXqimVlU3Dda1+mtgI5h+7S93zMGU03
fUuAAg1cRdTXvze7/6OWiCxFkgTV1HdKZHaVWXUJ95erfQISewQ85w+No6v7T+KPXCw+MIjZvI1I
K+OAKZN0ZxnTWUftsUcRDuAwLmRduvp+fu1exUTJGsMslkIDqGzqG9Ya0LJwGDTtttMFVt0mL1il
gdURpF7jlt8bRY7EoaPzuChe/m+dgImwxB/jXivaA0ZC+fhSnhOmBvkXdTQHHT1SuiRNFkrqNABd
IFyaKrmQyuSHCpPW9h29VDEF/ueb/UeKdoV8/1+7YA3y/PhGKqB34202YFkeu58xcqIzIyY90GyJ
c5NmvGLw3ZvfHHApJUfmO/yQDHZuHDqu1FUW6253fa+gyV+3a876LQnjSPP2EjtStCUqt+z5EjYH
rKlUI0AJsNXBZYFmiNcshxtXUqecFnPDbr7hpVyEUXQWcbCk/M6ZM47O9ue1h9spjZ7LCsvhzeCv
ixwPUasoNsRpGERky4h+vvQ03in0q8W0NTDB7BsSpKT4hy1ZoruFof0z/580sSL5JTGkXqOhRn8p
YYAmCwbOdeARNxwhoPieYddkw3lWAlhIW1o7xxfRUwzQqOcxTbCR9Vg6Y0rCLi9TRnv9D3hRhHs1
Uz9jht5uETuLhLxg+hNrgMIWRCqOwK91MTF/sEE+aVeDSfdJZ0KCce3CAsv6XcF0p2zGvXXao23t
hyPuCWhr9p7QISKKxwYXyq8sPNTqUhL/hmSzeMi4gfpgbyBk79MqL7mnt7xi537lQdd0JS+BfAgN
80YrmZCeZgw4i6tH/fdBn61MtTF0k+xyR+HRnJ/aJhB4BukfIrIdd1AjcJv2xJ7C+tmCBizlB4lJ
4K7DkY4X19gfiQgPjB0ze9fAgGM1mXtpdKNkQwuZZEZNxcRmYNnQbh5i2B2xLMBGiTgzs5ZBf/SN
Tyd3G+SZxmb20kXd2oLfSaAJgeugILsXC8OprLV81lVNqc3IeI0pSvdLMyQrxodd5bHvEHkruCe/
pHcPD37AT9pKlLg2igeLKwPdLon/AYOMTL7TEXC1sKtPxWRHJKIJBnoeSpWyEmfaVFkqB3DypTys
Dc0rcn5pTX5EdiTNTmFfq7Jc0jQU+4dyTdms8dF/o+/n2D6r5qemeycsXCSvrqlesQDUeIx9OvX6
oWwP9Bmkx8Y2XPJD3enlef7AehK07906TkryDiDzHYmaFnoetZEd7kzNCiDAbwnizqcAvj81h4TJ
JuQZtvOuPxi3wOokBN6Nm9WD3FbPocJ/vwCyRx4c+tfHCjyoDINAFk7aPHw7t67XMVKdoRyL8FLX
JI8P7CXSGu68gtI722EGNb6o/M4vw7Zx++xEFIS8ewmhFYEXYi6+HNDmyoJVk0SjhTUXtRhw2kIG
pI9fmQxxFHmx87wySGif1Bwe0bRwWRT8PnlO/GsKwzsLjbc5KV4TKtgS+vl2l7fsZV7bhi0TSfp2
QZL483QnH8XPHrwV+321Kaj7eqLmX6+3qwX/5s18b1iWZxMSMx4cIzJLMuPKlATGchDBwV3llacx
2rK7nHkl7V3H8hy+i7VuWX1oNe+Ra7mAyz2Xqi+qs9vUjJiAghOqoNl6+tRJq3vGMAxyScQY3AS0
WWrGNxRXr928yL8uW+MP6Z5VaCzvbNmUWBmOgcdz4j9gO3Hk56dlfdMc8p2ZrsPKZ8FXzaECUG1n
fDJ+CJbLc74BAIXgX7hz4yrueb7UqaFzPVzfBMVquRwtHxwMdgYMI6MsfxqT/3GELkj0N+jSXlSr
a/7g2SExZFlt/nqxjwq0ZYFIFNpMpPtJDo+LKNPHSmuLCvlQWnWzwcVTd3GS3xJ2Ltr4AbBGyq2s
D8umCDrBCuV3GwwwflXzBvU4fObXEmp5qPwWlsaVlnL+fAmlqAed1cb3dXnA55jWSAmPX4VzY+br
HZnuvkScn7GmFbStTh2ayWwU13CykjZG/EQ3NP3Y7z7PadurgMvQ+OZ+p7fS/91xsazb/MBVuooo
vy6o88OZC1bctjP04mBv973mS0vRuW29GCqh8HM+zrVYh8N++bkpTrstm3Mb/Kb1Z4S6kmAz/Zsr
LY/fK5V6nLaFmaBxhVOXaqayCYgx/8b2KX40egbr+o8D/ZtYn/1zZR9OwJiBuK9chNlQvv6pNT1n
CMSVyrsan4m3HoNA9jwPLhY0FrgrkP2jCpZ1N/9mfpab+RfoE2TVhGfiUuJ2mf76i4QT2bYUrZGz
u0rSyz18oScCh4VOhVgiUxSheqRZvV+TrTZa0WJIdnIrAK7Hp+CGRtpdbWyd0owItbN2XvPXnpU/
rToVsjTqZiR0X/WcSChzuaIA02cHqA9CdWXzjF+zosXhBkHbqSPFESi+J8WNf0tWC1YGbgQbef4Y
p5QX+I8KO9ApDrCX8k9ct3wXge2P8OUhAjujWnjKKPhifzHebFqmt7OvyzQU3i/Ld0On/8ZamBpo
YnjCNj7W1+qiD5kjeiT16RILE38yD2u4WDSuc8zaq9rpROyjC0482V5ALSy8YzSglf7m4nHgOai3
RMaPb3LAIzxAZqOVBjAWzUqKZYjzeEWTc4qfmQz+/o7XbqmYckfnMEFvHJw77zpitn53WvlhGJ/v
FYRFQ5s43TfyoGd/KD8+kqaVA7xEG3r7tADvpuBS7Nh29RhEBXXXQ3mLkQRFtTNsueUwY7EDnJlh
JTFaqdUIV4O+0lrHRwTY/oYgUTcUVXM5A7iOQdAXWfu8lEaITrKVWaqXMrXZx+3X6ey9CL+Nk4eV
LpvyxCDwXdkagLm0Dk8zBxGJaDdtODFZ7o+e+S/x5RcmSpKo+Js0WZP1eorf5V6XKbCghX01KKZl
snVU1j1AX0XPHox9OC72fOqURCFKx1F1IfUvF1i0vu0rTfxZO8X7EWePwhVE/ZCxt4VkUhy1JCZI
NS9x/SPAeT/7f/xUEPbC3BbjGl9crP9fJiQELAWDI0gWCEn98euS0OkeUc4ckj/yR3aLVHXWexuj
0nYQb1o+ENZKwPXResS6WQ7DwUMIa1JAbrT0Y7tn1NYu13awi8k1oAFFI9UoVP38XcMbm0jZUMoj
06NDB/sChe4eGAga5noOhJdCPfWji0jpBWQYArYlrw4mNU2Z0s5yV3pkNZN5gY2IOW5FgtCD+BiE
s00HZKstAupqEhdOFIWwGDRQz6qDO87y2AIg+nn/nUi2PC4M9dTXOQa3LH3LZopXIxYf2wr4ps0P
wQEomBD7oCWxzJcHvUOsHCoyvqhQaSZLXqpRy6EgLDb786Hhip9UIxQ/jqeXRjUG0s/GpuK80s2i
SFj+lSM9Barl56At7RLA4TlyDMzsGEkqpuCUqfZUeJLuOLOz/UjgntbxhSFhfjUUh+MzN1OuMvgZ
MbTpFzfBQS5zSEiq6hwYAhkPRdzAQRQgc+LA2fWFLasKiGzfeehOKdZx8A5bfa5b78H1fZ6QkuB7
LzPLLGPhJaoMLSh8yHZA32L48bQAUF+siYDsnTcvrDXO9ku5K7hk6OesLANPMAiZJa+UHTWNiAxD
dXxTkAAbFLaQQQT5Y28ojqyrjpWJUNSfg997uNow/5EU6fggw0bMZ8RkEjqt+xW0u1+MjqtcHYXp
vsfLuM6HCuJ8GwUWJqHrHaZjcB65ywseGIVeZRl1JvJzR/Mlw6kCL5a43ZX3JKRbClVevh+52pqY
ivHiUuypfSRAoet1WyhMC8GKbP5sO/9DMTKdW6rgr7+KOstXFGqqmhlI0hsrkb7whkbqqQUOC3gi
tPl6XUhaJeRZsCHwf/mlkHYiZVpmPMzNclOogEXEJYlgjcordSuokIxivIuo8qKLir3aonXc2SXi
RWpDHFhUGiCj30y0YHJiaDHaYgdgiFP505OCBaWAbeERurR1BMLD1JyIlBUSJLxMQmQ7biZBvD4Q
RB54Ku87718KM0fsrrDef+kAUAWFHFtbBpuh+ye0+VE0IPeb9ZOwgNemhRHmTcsEn+zAGRhdKH8k
NBNx5WAbzA8gqa9N4qXs6d1UkUP0ynwWmO47r7Zw3pj5hK9HgGRG3BRsfZ0F6NC3HVb1aJDzpWwH
w9jEP/nRwT88/ABVw0U4RxfmAfN9LUyH/vneK+tbZxPpClw78drR05DBgV8hrgVtrOkR5VJ2fJgf
joUvLR6T9aLHXSwMjL1A5RM+HVP6Yrg6LqSPhQvRaO0mZdkYCcqt0x6w7ePSvhZvtzv57LviEE60
1DzjlTbt+v/Su/PIZDXUO21ztGklcJf40OLg7yBVfEBQQrvJoJRDutCkYVg+7CJibAX1nK/l8rEw
k7rxWtc7O3BDasiEJwxd/rFq8GJPH05g4TVV4vdEkr/XPvcFkKItrhRHm61UEbuYcBsriROZLu+A
PR9GNN48dvPzYLjvI4IXMkpGRLoB4AWaZF/hkSTNIjFJ09ehLDad5f8uLofcN0amaH537YmqmrCp
qa7D3DBu70VyK1f+QFicXFpfkFK+kg7olWowErwv/eQHo/IzoU/bOjo3d0K/TXFsLu6bPmbj9HVw
bdwzv87JWrQfiiUlnLyThdO9bgSgYoIlOrQ/0tTLWVkt7AIGEQwSh26wLQFGruapgGeLNh7XwwFe
aWCwRQuXbVJdZRlgjfNwqR/ZJeGe+/vvE8iRRVAhQJLMRMTlp7KOzAYZu0bfGj7eJf0uLlqfWTek
ppGs2Ga5H3gLEA2hqf9mcawJjztvOTRTgscUFlzANCBoM9EtByJBL06C0PoKxdtVCMXW/6yvIVHE
RHIwtB2kL1HxlKOS51Z1XfvSPBCSq+c00OotYV0c7XgniYna76/uporVH7lMvvTycCXkZPsfiM7f
Z+oz+A2r6NU7IM10C/CONp08CKOGAeF12eUVdarTm8Zk4voGjXrQtzZJAu3eiFmAtsZD3fFZTFti
H7b+bI/qQIFrO8b8sWcaVthZzgMhSPYlk3WNPt+a1YxyMIMpMw31ylaLkw2IUXQw+ipNdylSK7EI
6cr+XaR47qDExD6gkpDFLzIWG7PN1STTjxr7QDPY5yNEvVSKT2LwrrsxHv/cfpI6UmAuE3RM3kA6
mRiXpiMYUTMHk0GsxJUt2yYqzEX7i2KRijT/M0TRrL1ADZkyLhWyhoUyUE6ZyH5xywsnRBsQnABN
HPSGDi3MdsJFivWJC3TaMs4cJxJDmCf+3cZEz+WqKdG276n89lxegflS84LfaFmKQ18a1S6EZapL
bTfzArS+DWCkKOUmD8gUo+ygUfRrHBTsTqZeVQA0yY2Yj1iiuMiImpwS3mBQbyPHn4K1Ey7s2AAz
Ipq+NiRtLs/xZNRx/jAv9dAi9a6VpqOpukuFHIhQvJF9Qu7LPsyN3BgsPWTShidMZzscztDP7yE8
J/xtYPOBUi7oHMf7uk/+v4ZOFPbLT5lvlTJ13URTUC3l+ur2FLCDu/CSJ6QK9jTTFxdZPV6sJkLA
8sKh0dIkrHUh9M6O6T8KNefCW3gFlTwfhKdmAsmJh5p+JszJR2Ib1CbFbLhmh0GbavMRul9/8YBw
mP7Ab16R0J7FsXfPV8OxnGm7YIUz7D9n8h+K6Wc1mLJNevr409sFx+Rx5WytOJ6PvCIM8DJ542K+
iH0qPt9+vj45UDcEDBIkOooe70CF+EJDDpncWHsXi78hpW3inQ+08L6Dt2GxOTPy+ZkbAjqFwajB
VFfUJb75yXvInQpUdI2lBsRlkp5aQpBu75GqNOJKDJrMYly+CFIFsxV69hjbf2kqi2E7I/wrHhRt
YHNKyxSu+Ei0zISy1BF+LCjqDNWafhPF7s3tzrre2Iu5QGikPo7oBgmAnbm1Hls83uE60fgpa6bJ
BnnGetixeP3V3dGb3t+847BTDhJOxjZB3P41PzXRvLy7wBqwe6WPRtJyRCre6oJxWGWzrJ6DlBy0
Yz5QQd7bdJmSA+U4YZoefB68Y5Lf1mZ3fa4nfya+t0n+VBC27ev/3AfHvSU7PqZiEHHB1Ykno/Y2
apMMXxKrscDgTTrEBowDGKjhPvr6IzXp6BDOawJ6sdt4lQSCLnzWFErLcfgDgJGV8h9mNGqBXH4/
ccueGXtrAGsW6ft53cYWkc5witFvNU1q97gLSuKSv65O2ASBNodAy/Ye6dm9TyZ5KT4b436aDco6
+od7PkagzYlktG3JCVYQ6vSLW8bVoW2EXCuKecROkPYXz3cBfqxy0avwqipBF7beA42AeM6jmXXr
/UKvsq9NKALERXmqTpsUHKczyYbTr+JXuXq2q6pNch+i12xr+g9hs2MeIAAwfY5bsYQtctgmHLpT
ZPvHp+u48C9fn7A2OdoclrG/97XxxM86YkyFyOclSrGdEb7xWEZiFUrLbkOhTZjQBOFnlf1gelwZ
dTeyQ234RYYzVTJIkIlkp+HS+v20IHOYYs1Nc1n2688PC4z+VvGof9cXFLtPfjc3v5J9wq5RD1Iw
IbJFXAqTqNObNQU+MbbWSG4tM3k9Pld/E94hD+OaM4r5AaKj9NZFQNC3WhVhPKD0j7A5VQWhiNj6
7yBNxm7aWOiklr/n22DlZQmannSsmZgxzYIcIAvfO9rviAT7FPXAnXdQ1q1ijNILirJULyhUEEwm
zgN1rJuvpBdg1RPftavz/ni6WZd5FpYlrQyiqect3DeBptSdVrVbBE0xWRgvhrg6FluoEO1vhV0Q
l5OL7ZkhfCZ9TaxPfou7tnc5QPz+Lxm8/HS29L4I9+tmnDGQmdrjSHnFDe8dpZOQAE0PYXtj4LV4
hfz/OeU7jiYTRO9nW9wsTCNxYPnLwkhRk2wK93SNP3ZeWjwmGFV0DINCuD3tH4pnIs2RZW/prr3w
jtLgRv738bYe8/Wu6NVU7N0IVXSUJQujH8o3atw/6idplPJi/HzWvfwbnxNI3regONb2GrVqcn3j
lpAGK121IxVYRd/SFwY9gk4w4lZi9K0PR1gJlliwAWFTOG0a4X9aZetYXk6sSCA+PgUEXSMt60bk
oulGxL112cYHiTsPcJal/Za6OcHBSQWhvHnRRNAaDNVfAZIPzu9tJga1BDieh6cVC4MEhhuKekNN
O9FYw4mPL86b1RzOVTi1BjaplzYbtu6bHPv1ND5wyYOxl8L6yk0lU199cTYTpO611tiZapFFZkBz
RbHu75xjcz15LTYvF15knur4z41O1TBr9QuqQBeSBXDIUitbLr85/1tOHoRDvTFh4AeuU42pTg4f
JQYzoZXjieLH2pTh1YsBydmtaGgLnrtOxITU2jPTWbQ2p5pTKtLuheJifl8L+HCPBM9YsbEbbons
7Sf6yYE2bT4E3vdELgpzZZNQwwjKtThYHMgE0bRJSeFe8vuIhAvVam8uKDJGQOjwY6tcvVx8XSaC
xFbo5h7l8p+EyDwNRQhU9JzJXdt38/b1BvnRxSZH3kXv0LrWYkwTr1PXinIXJlTz9DsZboSByxAR
PWNYMAUx3Daql1zA6jCyURKibXzQdhEImDmz2uZ/N7b2HPeNYGWStpfyge+LdhLTDp8z2dBjdJpr
7I78PeclaH4KgsZYE45yApRD5zxmH5QFAt5gr7WQY/lYIIPJNZVlUKgmuCBdjqcUl0gR+bDeSP5R
cnbKCacDoJm3rWZxZHuJFq11PDHkhREtWf+BGsuXr0xGGwDhDucOkSsueb252bliEjGuhjCDh93O
NNG7Td+mfDtD1BoW/t4kcTGSFMC3zDSLT4cuYEqfvcnWY4DQlKHJbuqG/zmhwUg1e9dMA1UlqUwr
ZpM79AQ+6muvp9jEV0JSKs83a9N2Sk4MIWaYZe3bOPKVk62N2R4fHJM7bVgSm7zM1r+4zrRWP4vC
d88UQ/XsHMNLmWxzrGra8ZtRgGUxV5GPHMXlTM8EgbUDh7xvYs2UeCYSUD4dBMH/PUH/q0/rhlhj
bNr2FDqGUKDUzzZsWQYpIq32ZlgOqQc+gaagJidVqQEqIgr/vqEXKqlhqhXUjs3J+IXuUyPgaKoP
lPKa7SLIkXdXXek1qFK1SChkoQHa8s156esdl2bpM54P6+Cdhz9raQvCFHL66xN/rR9xlIqcyhnU
hVN7wLkZ9ojfCVlpm8vMk/VRtr9VseGKGh6UsnkZ3EeXfLbylgTFT8No2SU9RTddkrXDQhDkQWry
gzsZh0lz0fXPsewMeY3xMtNSYlAwO9XxEE4XkmfpuVWDsSy1NFupoOVdM0/dPl+j/gdJUfBk8HFe
JrLib3ka1kHi8cmMhVYM6EPMODAsdNmKwvSwBruTfzjePqVEGQBzVaDCOArOPEExs+M6vBBVIZl2
tVeCnjRaOZncKs3GI+YMKmryNSuE9St/cIKn+bl9uVpcH6mfam4D0SuY0VwshcVEe7Lhl+Kbvg2f
jxItHoTdVUMBeLMGgOjby0if0VEzcl7qr4R3kn0nfflJOWdjZ+myXk+GmddA6VfQo94kecYkEe+l
J5atMzF70gHzSBJ6He8eSvU4PK7JhP+QGz10TERPQt4ARE/sN9SEyvZiFWRdKS6dmv4UeHrNxPFD
rlc1USBQQJHxSoa2WKOunt/dUBZs5+6YN739UzpR1slFws5AhmH9rQ3cL5gU0IOPnq3QEsCf4dMY
LxIX7mjicU/kSR3GU9jFKhm5wkYUS49iZgz7naNe974UVqulAK1+ZxgzjOj1t68yBFl78gOdui4b
qqV1ldgpau0JAvrlml6d7rmzlzMIEffknK0PIAM78FjDwdJzo9AfiMoxz5LXcZuplW70rAU7bwFu
xNCDhgwAI3DedNsxEHTm9J2wChPfxTqnPFAuYAoV/i5UsLlBDl4SvWOt6SdoDVL9jx4wHc/l06qn
O9lphMzEj548ZpAuIUiW9h3G/j2V2AXWu/G2tAqIKBHMH7+6hwjsoDTk/gbikBumUw98y8NGrJMt
/5vH2XZfymGlO1G6gwaolXMY4gDVwAHelNPNWALXdf99SUf8HLAu6nxKFle8Y8xM3tsSOUMSuxDi
U/19T5J1MUM7GiSouOfkRlJoU4bd93VqFn43MqcYaqGIOZI6jYIm3/yr5nYtmfOwG5Rg3naiS3Eh
wSLXYd3g/e8bSUCCVZE2IIWPtgISbiboxfLBcIWiBedcURO2vCDRf2r1pvNq7lYn9uenYh1v9z1k
QKDkgi68tr1tkeTBI7RwCOyU3pE0oknAAcPTIii7+qs/ZBMbBUuGZ5qalQ90cTaQUQfc/wPg3nRZ
Etg2R62G9XQkNW9Qc3uYHtaEampOeDS0cK1fxuT3AJjxJmDkKz8ad1uj333KrDlLDP2HIdfo4ECJ
vnRuLQoDBEpqc/LzOv6M4S3tUx5i5svXcWAXQnWSshXggTBOgi7dCn9SBqfPn2KECCzN9PgqeVHS
PS8FeAMcezdTNChUVubBl1s6BZ2RSSGCw8+t+D7MzxNbD9HRVULMaOP/NGgap5YTSnQYJ3Bz72s7
9gq57KkwitG/YzDGMVWWApP8AOWRMXmvwRAj6jq19tuMPBPJJ4QLAL6nPQD5jGTL3DmPy3+oFcWs
Zxve01uN0BUaJgkLktbY+55RT4CPzdI/tKqNaTc4lGY1J/MSknjzTQeK9sh5Yt6z4u9t2sAwnc7Z
FxHN7hRjWt9ymho813/FVPhXFz7uHGNPDrNXUCsrnX4qQuteYKzvXwgolppyBvDzHHUVBAGWPPgE
TDHkN/bJv0ctoYAh0TABagn57ABxi+J7jrO244V/hV1o/ez+7z1bqYOkwQ+qauxyYv4f9mz7Qd8K
/TEZchonOb/L0+MiXF98X9jWx3HOH7+H21hDCBXSjr8fybdbodMWusqehl2vq974W02WxQREJx04
7qxKaa7d3HdQqvChmiEq2ePO+nkqkz9jrtbCkflgfCa1NzRRI54G5ST+XOUgUYLFoBvI5bgrIKJB
CDq77MwO/0DURLjv7BZKQY8OO5rbWDfUGCzHk3wngsZr+GL4XwsF8b8sDEFHn1ICVsE6LmMf6+vo
X+KlQOtzhQFG2RjWIomvACAgHhTKQfvHh3vGecO7KCH21pHooF6A8FTkmovCQparoKCqxJ1q91BW
ACmVXNJYoGu6LzAEfMJs8ETFss4ekDxn4EC/tOFeq8mv0YOjr1UIMqQKE9DR2M9qPHkKnnWB04hB
OoYzpMHIqdu8LafQM5WBAopLglFK4tdJP2y0XhdtWn55vk0UJPT8zP01qjEzaJl/HcQ7xw464xzc
SZ6ZMODqJXpioJ7ZUo9WJCBh7OLGHl/3w+nxeFtIs5PEQQyWrC2ToF57zbM0VAYyHxzJ5sDf7A/g
gWqHxqEOO9mvt6KWo+MDlADydkAuyrhw25+AV6W3L2xJsj4B6dlKwJjJzye/PmDrv4nYvLVYsCDs
DDv+y9b+ho3HBeR4HkWEXMiBtJQc37Ay6JLH/r/eHOdz7fmvT5gXoDz90s4Eca4X0P/Wpa8pZOYn
6iAjeOV2Ae1MbEYSRABWUq41k7dPrT1NcCw+88M8PKBUXHvYgI7a0Ez1HhlEHU/y42c7m9+qC+VR
tgU1UV0SYS06A6RaqK7IU0dU0vmi5GKBTl2mzzKlHsyxjWijCOoN6LbmT2cOQi5XqA/q31CW3mdT
GcGwRP4qZct84RQMZsrk2Sy0t8pbEMPz5IbXQyivqPLWyaicdM7mzmJn6BJS7PlGtvlSFFDsYIL3
VAbxyZ0jXcJlCjPKGQ9LXjSNICViuzMgtWL8OGhrcL0MyY0YR5s8kRogTVpzINjOKLrC1r6enL23
FC9pzGai5cMWuxoLWY4h9ywZo4vLbzmCJ1FexzKB6OF6LzmgfbUidPmnK5kdzeEXXlapqcZptOYZ
ZltBjI9wylQmROPGlQgfxhzr/eWWvMKmxu75KbIbLm3MuHOPbTUNMF0qkgPBMC7sS0WxBFaEGqxB
XJcmx2tITGvAfGy6/7vvhre9BqVDkO3R9ykhGqIsMAg1e8oo5UyUuOvqZmyPE7JA5hnsscgnJl6v
eVUfXb+M/+fwzFsJXByYNA+Ncm3IYqFgjTR+O2BZY54NutLX3Bep9pW/xwjkCR21XJ0hnoStsAsX
z1uVdISPbhot1DkeoqdJWzf/LPutChkDjp/ET7h+8dGBTqhdiYj9ASGotmbm9ZdsV33sAp0m+0mL
ExAJoYEm1wFuk+IC558uDeypTfDdRSJic+wTUBPET3yZX/sfLU1Dpren6WT935oivPRn0g8o2r9Q
+Scmd1g73akY+YJsRv+5IE96BaFNRyJq+OI3TZVZbel88qGTyetca2iVCdRNGSo/sAHMsYKHK+To
Zj+9hOIVXGSNRkea/8t+f++jk2tmtEvr6FkUe6pwp/TAvYc1wqoRaRyyzHUFHOzLDs9eT7XGchZz
RsfZYNNTIKPRzLKnYG/6HN0PCS5GRpYWRlKVl/OjAABOSug2P/qkUCLkRwVc+Y/JjMpbrD1uaAqX
+mb5mwmMCe/4JdvRiKGnMQqdkezN/j3aXGz5Z10l0gWPKW5uRhPvGcAqhjrCZEkvQF5gBWMFQz7Y
cXD6Pp0B23NxEcHVKMCCzkKXKRQY2yg6EPzIp5D4y1V7tqnfX+KEi3yp5NiUEKuxLAEVcMDxn79x
+cE9dVXriyslbKkl41LoerXUtZpWqA4gNVfZIbRfCA3sjBLcXwicnYET5rxY8vkvmoJqQ9rL3Dfj
ArgexnugvlywjbJuXgThTUx+b7+lr5+a15L/QC1izS6qHPktkuT3SMyzoB42T87RYS6mx55dyRqS
sAz+fP/+y0tjpX7PvvQ16M19qi0wEoUKauN5WUUVTY+JSuC1uRO36acWvS1/I3be/OdTf6RaaB6Q
JDZpPyPApu8IHtIISE3WoUZ+ik8mhIv/nFFd16v2LQHHINpLBoIegfJPaxdjzvlwJ6TfkQMHihFv
Qprh7YRmzLui09ewTCqDZfCAPWyiol+QmDCXclinS2m8wpIOo1N5tZHLsSJXL8UkoLvZE/7+oJgK
az5wt0hHnyx4dMVCfj+/afEozoNu3tzPGqXvPPxa4mMuFGS7ZXRmhtlQdoRNr/3iW550NKdLpIq5
e34A9TbtFBgbdlVrCoP5+qGSTuhjhPUF63S+Y1XqhZycvIIjX4cpcPOOqLikBGaC7WYmueJssOoB
TxHa1t6od81eLCCOyA0fFHuu1MENbvk0X6hEIaugRP+ul7fSVCfrsBTw4Xa3OrxMW7N06yLpDsk5
7LF+VjEmO7Ooz40s2WQDQ8JNTU7wKTvm09iyEP39Z9II91Ff6WPGGBsAiM2+DouSNntlyCJtMMyw
3gqOMh0zI9+IsQjobJ+7uJ6xkTa3tm1XtUJbWHT/CcvPm9ySMdzRaXbSwpjQjp5NrGb+Z3dd4X5K
rKpWKnneT3JRXqolyKrVHcCmXf+puw2YFW4x0UGWiejxjODJkH/+6phhwXOQIPvGzZ5c94gPmc+8
TfOlHkdTZjYtVb6TTILTs66TgpC22Yo2fZM5CrD1Wq3dxsa/AQUbVh2jPSHbTtXjpy7IKhl04arr
cRqOAZyrr28n0Kx6ls4a1EkhEcVPQ3UcfBL2g+cWVcZmVV5ni0TJFHyo4GVRe0IYr8MUop+SVznY
fMei8JI7q9c8YY2ypf7k00M/Ot1rdOGn6f4vnsZy2N1/GhvLLRxuhZbe/ibDv5T0ULraVKsEXiDT
AE1hCLj+WcZyp2eERAHVtHfVsfiHTOXvRg3udCIXq/XuAUm1NSP9KRbncGTmvpfNamix3W4VjLyy
tHM3FRpMfvJMt9O5Ek9Mppy8O+FoKJ6ShJuEGZ/C7YQJbqDYPsqMnv/CQzDfk52LZ6TOwsjQJpPN
KZfWIuNxCz1nKwI4OLnftgc5Giz/KkJBkh/IPW6nXDr5GsNF2Fj6KCk20PiwcxBTTK+zULMJkkHj
WAhgHf/IEP+iXL9BGBvwizcybaek15LfjR1RS8VEvducKOCg8tK3H3EBz/DcbPayko+kxmBxmN4B
E7aFcYUiUWbHq8+v2T34/WIvXn2Ujhs4uaf2wEkal35K7leAdLPJl4YjcSq0XGgGZt3vaGoWEnpX
4ylslLVnP4qwjX5dpqMwTUsj+vNJQpjriG6zhaL/Jy+tfDwQZzDVVaTIrnaCSYlINIeYcGEWGVir
ONTnQv897I8QTzOsnEFhZ5iZOTDr6hkGGhqtsASwf429OjtMniF/YzTHRf+aft18jj8/Zyurabh+
YwEgQ0IQ4us8VNthCCupFwFBZZjXmQxXNuarshhoOkIUQan0K2Ux/cTwcJfMZEAT2qZMAMToSsGI
Qbg3d1e1ANKtGZteGzhS8MnNTmVOjmtikaeSNcHevup2uKNFEK17+RRPSjNzF4hkF6PO9VJ0gOKf
8oBaDtq1BE6pBUXjdNFlUZTE5vYXJdpRhGA2OUwQgh5bY1qWVaC1XUnHHWmlrOoeWLs06xWxflTC
6/Ma5p5ZVhKj2Phvoy3Jeuqx25iCPaQxu31xaFxTwhE+dmL05UNDLlkqoD2erS64T877ALsgwqgH
Cq7ssaZsIaEqYiN5/ZxMHC/j+eRGHZT8UP9LTpafci2DTx0YedNQa91/eWFuptgRnktB5aPrizO3
4qXjPjrzIMKLvqWYb5k16jPeFSz89HGTMXH6vuFo3wPh3ekF9v6pQG4gd5gQZFKQI918nDWf+GgN
P1bKQsifNMvX7xmU05e4sjLdYLqDS1tFl1/prol+Zoqc2hyFzOg51gG9WKjs8uJedCx+0TPSa23S
Ee6O9uUVfACNi8XLXbYkgjllDuAQ+eBocWZRwZ+oK3s8X1mgPgg26jh7r1mLWNZvTWjhXG/aK9RC
bRduHRPPLRY3IM/syi3a+7kRXe/OmCr393oxizKUd9vhw3qG+dEF0VpJXgg9F5utzrMaNE+P+k2A
/mQwCuVS5tm7tXh2rooJkaPYEn1chXrsUX9KllGDwqJZq/OYakQQMTzVbrUt3JcdglxzGGzAJ4q7
PniJIRTonFDGEZc3Plhc6nb21xYo9TU9t550C7TdSlDIoF2itUxLNNVGUKaDM6lg+MubYQsd5GCK
RV9zlRRJmKelk85mCEnx8MfnOHHKfJDu0HCQiO6RDZen7+KaZnUEQvrybULhHVwQ31Q3bq5nealE
u97e/+optrMcVJO32YmY8sJDqNJ5rzVqV/ld0gLcsnHivtjqYMFGRnR0WFu2t9kimERwr9pB6NuW
O1t5IoEd+Gfbv+YEV7+tL1GP4e4ZcoPbE7RqsQVb47Z+ecOHqateIrtCr3U2jkHtMB2Cmms/x2XI
5MSd6SH51BPVEhuS7n/QciFI6MIKI5G+0nPwACxuclsw4vj9hSLQxSimzXy26rwkIbRW2BLSRH2D
SmGIa12juyCk+wHuA/Iw/TmIMnY23lNaGWCsUg7CNIUaeiRycnLOBRr2z+3OyEpBeGl9BoHjWl/G
mUumgt5eV9PWDvQZHC5eXyNxCJZjbg/5w4r8eBWNpzbqevKSf0dhUTLNjcJUU7DaYDm1xGBljG02
1a7PPwcu5VeldKcLEK5VpfJdSZFakygGI1FN0HeFlm5pIrEEMDrHIYXoZYnIDbW/i7OenMNPWa3H
CdZS71rsLG1esXijRizcR78nLi8MjQrRGEFcCQ0DuiOGFXwaBQ5QguSv4no6Po6BH9kS1C39WcOu
bRnJKWXO0yoRLHT9y4W9pgHZzUv/W1YMLE3aukLnWeF4L2dcTrD5KsZLJFzJaNMm+KaQ4874TxuK
vLY6sSv4ty5XZ1fBseKyjhgfRk7r9WsTXgVkHBboEpyLvXpgmwCiZZ1sd0U/ptBB832GiR3vLxWV
HY/8xip1XXAw+Lfxov6i908BPpVVTwB3dEjij4EbPmzFnUmk3ZnBInAwi6aGZjj0EIdTOiZaBXcB
jLiNES6rgmYMSCZQ4ClGusdw5iTcpZ7vmChtRIR0ZUGLTyH1oLAWxK7LRMMkGLkrhOPAVAuhkK6n
5aXInT0v8ShaB/ZYDzzS/6nRpQ7BZhvt8AiP6Oil0UpxSS0fdFYU1az2yDUt1dm4skCAx9Xaxrty
keGUQq7+k/ZSV0tsqU3L/bda7ghuSTnhgD9au9z7KMLITYzpoQZ0LHZlBEFf38w7bYTSXtqBXzna
E4xr4NqGKWRGoW9muygbaqhyJNJinHTVcXwBq2FHR/qJM55nz9SBt8J4LMgVUpTGQXrmktd0RFD0
PoqASVvD/5SS48wmkkdpxTbNobCxXGwUOCi/BShzT1+jSqtPtQj4/kEWWTXBq0ROIhEb1IOMiHuN
Mi8Hk13+l2XBs7iUWWcwFGTLQ2oRbkfE3vyxdNXagK+S327b3nd+TGV4r/PSEQp2X5DYA2PxeyU9
6/NnnZIpZs4L/GYkaR9XdH2RdU9cUtKQfR5RM1S2arKTfwDdAZ6XKMgsB7vX86VNbWjtn0V+fKVa
CjkvJjTI0NxWuzLb7Lj4FyGgWnHGaTRL2gQwQDCz7GuL1WEyFny2CZZ6rvXMX8uWS/nMwfiSnBDU
bJzl11f9/gT8XtDqC3ZJpkoK32YDJ8/jU6H6g1DVliNCY+fdSjer0QTXQGxSoo7dfbtpDeAtAkPt
vuR1LBpcmjYETPjlC5U4uT8LBZe9H7PbezrcX6lx6J8Tnly6pgmznzpoZbiSRLuGy0Lc87WK5ncW
xnpySRD5kb+AnKA4WNyDTuIps7nH2+7xY4VT5OizCBJK5/KEoO7+dWSk/F/0bVWhczJhwvOgo4Bv
9RV1hQOv02dQoffRDT/OrjVO5fo3TTcolUfDN/qQrDHBtXmkFimRIg9LSXcSYUQB8FsVNbJ0R7sw
uYTPHHhy5lDOSBJvXzoQ5u94VzH1HbRPGq71sw/YJemodSxXoCSNOvy11HBF4p3DRew4t9PBAyvc
Zat9VQNQwqLhZzwjnoWbxS3Nft/b7QA5O8lnPJne3467CAZ7i6st0l6GeWyqUlVv8yi8SWlfhLwt
O+iQ6mHb9Lq0tRM3tM/Qy3Ia3T/ORTA0cif9rmEeVI+kFQsBs9y6VqMN+GuCbi3dk3vtqJZpDJbI
XmGbcn0DyMrZXl7GIqQwlN40Fo9KbbYxKiPZERwH1E+Af9aWBvpa2MwttILiTCdE7pfa7DVzH/zW
HnmOIaPRnMUQyfvnbTurNV+I4HpaLuEWRw5uTNqI4XSUGpI1fvxe9novcho4NORu6Sy1iqRgewSL
qoz/zxZ2FkcSLdeycWsSrwE9n+lYeYtO8X9Ye4k8jd/Rh7DZsyx27HdAs+X0x1Wjyl9DTrkDQYwK
/XBWPBPWbqKZXGcAILSwwoxeStaL9EEaJDkd7toqflTaTLLZMpxYH3kSOpDfoadXBMtjT0J4VOUA
cf0ThoZzTWcZUYbEEaUzr6bV32tcG4pqpHG2MfLx5OQ0mDH31p74zBqkKoGF75jtir6/CCoEdWxj
cG6UPfMPDpBlXcEnWYUEejsUByUnNbKIMixTY3mc7NNctvFXJSUebtaUn2TqDolxqXOPF9AzqR7c
5SF7CSrlA6rXbtm+ycNrtqYxAQGMsHVsGNS4mVX5WCuhCGMVfQsqLtdHUgFa9tZJamMp0bMOooYP
+cN8g/kwbB+dePAJMbOtsGX0cAxW4ifWhaHx5VW/tMjiAzYo4zK4BaDwNF8zzwY3k4VJx6rRnmaG
NkOJDcGQNZ7vel4WKlw9gtajVKQUp9MLukVBY56k29Z+uI853GFlOLD3fNGetDWBCzrmU71Suvxk
ESx0irVSGrXDLwB/dqCdtcyNyqyq1TuAnx35dm90Vf69Nn/PCU8/iAETzjjLMSksnz6BVBDzGK3K
Alom9I5omwKC71Gtm7gWgHF8/Ls7uS8d4c9JWIjeee98fYZcGGAuSMRbYgfjaQgwW0Zb7V7+uGpr
aEigm/UTO5oGpnO/kbAv1filh/bC5cN98W/2WURWkZkYSTVb6oGgGKCtVnGucyOJLjK3CTubiAYx
DC+8mOEIIcdqSwKXmfMqi0jtZQI0mKA3d7udR8Ki0Et/iE4W3BfTEEuX//LEfgsA0FiP/2YawNk8
bLaneYALxxnF2zVdIMIe9uODp5ZXv22cTKKVgnDXZzqdZbYrP4HptcsNKoq4zGjoyovFVm5de3gY
aG0hl4PoxG5w3MCJOQE0obWvpPmBW/60zwTVlZmCRnttLhKd+xmzeeAtSYAm7tuNxogL22ro2BVY
Azn3S+K0qh8glBEHQFiq/yrv0eTDGiy1+EdU/CY2Kmfsoik7GGF72YBQekKYrm7PO9JzW0HIM24V
0U4pvWIpXBBcmrhKOvAqy8ci0cuUKysn0B5xMMOUOsWcxZvD0UaXD64SOaxc03fhRqeDAuFNNQYM
O7mPyg5n+Io80Cidb4GkyrRA7wqJtt5MRcDtHW6CNOZQjTQ/rWPIwZcZJe/btCfqG9OjVKmJ9GE6
4wsdwv051FlthY10k7Avl/6i5nqGKgfryRMQAYEiZmT7ZVHdLRLzGF7RlIlUvZuSVDeCiVS7pTNp
8z8W8WI6fjzqBtlQmHZRM8ZNFlaFA4C6B9uPyh/Hzq4laQhBggnvgIIFLpxPzlj2fxm+05TCI08E
NmnsgIswRZlZz8C4IwFpD3HBhq9bwCJbd4JCESFRRtlZB70Enw8jvNzou6s/N4hJParKt5Svf5og
ObLBqpizuTN69F8rfis+YX3cM1bUyc7s46AK/vh9lqVGq1bLEzwCS3nrXOdwkGf7xaeux48msoo5
4uS6XHuNfAuZ3p7q7rKdYmSzGPjUi5nHWhA4jm+ECGApjVQ+elOgce+t74TyMkuXe5iRPurtc95n
hW1LxYV7txo5v0OuKwwkeLvqG7sQk7AAB2uRoLyG2SVRik+zJlTHX+R15O5WuuCLikqzjEysNEJJ
2oKZFzqIfRp0EFg3dsLkZMvTbQp9UA0s4W9Y/d/cWLhZeQcsoftlE/JWU9cEiPd1nL1RpKBkDWgM
36CaR+Wx60LlN6xtsMXSxafAQXID+ahB0lqHdMvrfwXid8vi2amMWvzrGCilySiG00tN17Xv3eHx
pMU3EP60D9lbdsJTE4pZkii2D3lCvhlIC/ilcTGW6RiJWAo6IPKCMvff4tEWQ+OqP0aEOb7Xz1ff
NXrSaFn+ik2Tk0zjIyNRUArK6sqpKoN7QS2XLggjktk5s/Lf8CtHX37Lpf1o5RnD430bbZ6piYAN
Xp8gcpju8P8Og7dT+3VvTyZqcSwzN/Kea6+rm1sN3WQ9HkKIFELIZ67l5kYfn/pqD5j4i7nJXb5X
lSb9ViFKYet6a1dw4XEZF1k8wSOcDoUMZUQ208vbVzAhaR7GyQoHCc1wrAJyNin5xsusWZ6C6K4o
mjF8uJ/FDteGJULbmxuhvO2cwQIaIjyfDZyIZW5G/+hIM4CvnJBU8o6oynphiW6Oe/0ORoJgQstA
yTbdHgAxdvAU5IZpE5CQX5HOikpOn3jIY79RxJYsr+VTKzko16z1CaKc8gDdSWqG7CPcMA2NFMih
6Zrwv6zlVwB4aXKhY/o3l+0Ptp0pPerWJo2FEiKaSJpi3OHXRWQ9pj4KqoOJUd4v3Qr0c7XNwQac
b9OfV9/duicw9RkGUEhMZooV9TkJwZ7aeM1ZD07WYxd1Q4wratnD+4tu6GyP/KB/G03ugWYO6+Vy
NMvD60S03Kiyk5YvF71JAzzs4VzKA2UhNadVc7l5EISkbStVGELacBtemd4qFhIGCYo8WPlu7Mvd
H6qiFwlOVcaRz6HqnGqoCs6rdn0qx+Sc+vr/NJ027Lq6miuvG4E6dJsgktpFFH8Y7Zs7Xrij3XzO
275FLHpO67PjSOgXPEpAwccH8/dcbTVUrD5FvbEjkezmlHTsqhV9aIo71D/AruuXOz2ad05kCjOf
tbLAIIVsTADeDn2L/GqfYDqHN8qwgzn8XZPqvaUWHvtQRLSy26D2pEzKiEsEtR8yZEaINYNUySh8
ebL6jAp0tEJ1IrzcVk5ad2LQwEMpmW3145ZV/FcFnqmcCX8nPPlVD5cdBexnP1/OjS1OfN4Meo/F
TRysiX0voNIiJzCv0eEIJmXO5AUZaezrrxkgB61gk24uh0za5xnhtQGq1XfHuFyV4t2x92beUqls
mvnbrhq9sIcPL5XHfPE+6wpOVNwHIQ2UxCEu79Rw4zSey7cznevLWTTZglfFSIZzpspshnc1za8C
JhNa8jzescQ8pgc4T7chwUklesJ6K/hybCmnaeVEOeBWtewupcq+bTmasqQwJAh9uad4YC+SZvzg
JX0Mrg9l1LMXPbpaVCqZNExHDu0QyzjBZKBH/9HLhNJ6yue/NTlfpq9Ka7vAC9by8Qv7805DU1EJ
Qxfoig60HnRJFsJY9ZWLPLsIwLiVyzO44q/jJqaH8L8vqTENYmySrA7wyNG8TNFc0ahVQ6ZyA3ib
r4LY7sUrKDw+L6b4HJouNnzKay/2VuKEndBttH7Y9GUFWlr0528iVq+koDh7p0QdXcHL3acE/7CI
+5THZHBtvYDmMqA8ama97/HMxZ1xhcncz/M6N0klU7+lvTafYriAIuS1MCBQNkvW+dNcc8BkPO0Q
2HTW1/YRb34PtpmAQ+TfB3/AlhsYcXc2sKL/p1TKFlxkW/Lpj0ohhopIFJwPsGpE/hII5mEMpbZ2
u3bvcrtbrQ79tX+lNQ11ez5kxJsNnE4MqXhZDbUMb1RqVU77Aj3R4188S//OgwuUX4JhccFRLx/V
lTNuZqVqQAYhz6tuGj0TPEGbpxAXnCVLXOq622oTEl26Hj5XUcyJtT7sr5JY9BbdSvCuDyIsdJnL
o5aDpQADKg6Bn3P5SlFazcsxw3B9k8wrtWLFSdxKYexZmS4cpgWzrS/gknUySjg9n0WvUY9iGXnZ
eFyadyGx+zUyD8KtZBw75FkXxv2jWScjqBP9DaJJi8f2nVj2Khv3D4UN0WIXdLoK2ItgkvfwhZtK
7ZIIvGDapjAlXpS0KfBmENrWFtBNZBT/eU5QuUhhDNj0Wf8Glze/T60kfntnCWNykiOI3DkBG9Q+
9TzxyPqdVNAkO7wA22urJDN0p0YkHKtOI62/+1KFYFkoEfB9/w/TBBZefzx8ojEm3aHoxdp3Nr2G
a/E8lfY9yyI0anX091Pqfk27bJvWZInc5Jc7eeUcGGWWxRaKg3wYQa5aXVf4kIF1LAgKGB/IQmHw
5yyGhsBJf7K+ThzPZFn5UKcu7YdOCPr2dv8Zza3JjiIuDZrgqzBBzed1SUFn9O93jgZuBTgMJaJq
fIC+EuRbEoatCijuadsE+jm2rbjScRdI9Mft1fUPz6rLgMkx2mk0thhqRk63EDEUlKHtzg/c2XE2
h1JUoodZ1GARiQ5jLy6Z9XORUg/o52GTf/L+PkxO3/EfcPIxWujah5pOhUnyMdQXEv0EuHgXOG5M
lqF7NRiJ8j+rdLjZfbc5vo/WxYLgdpkBBmfBi25T/fAGdL+BQkhguybWD9qsT4zJADcMqk9a9xoo
Tf0bJDGLWtNlknzHh//RmC4DaqDeJtWdqZSuvQ7zRpHtGa5FjqkN9xJekmY9bnU6rVBtbJsQ4ZP2
bA32+2hkrA9Q3hmdlEjRdqpqK6CDs50D696PrG1/+754wp1RXb2NiTruf4AshX697NuyJrKhHfrV
UHWEirqMdqx4NCqkktCHf6zLfSilQYicL9ZLSEoJthHSTz8hVmVWuq5QcGzFTVUa/6c+Vv5LGOde
jsvHx0PPqmqF8MEDzu0crvJtEBcGDZYj1Q9WYiYo31HyWBG7D5i98kcZeR63pOubbETufZxCv0qu
7V+YYCjdqlpMMSB3hoxER7xoT8qkn4rYUIwfjhHB036quWGEdT88RE0EUys0XvY62y6nP8SNX2lN
LZml7HzohLmjWlTa+kdiGkNj6rdkjTMWYHD3GTm0XzdtjC27DRZP/ZZdzXrlDXOtYEVJbV3WDI0A
eXJH0UufEwaPARnO3lTkwzdTR/XKfImptmfp2mJcd9gj5YklrGRWrTEJmo3fWNVLHWFMvb8KDRO1
F1FNKot7vcbln6l5M6exHjrNdHCn8VZFm+0a7bhfi7KkxS6u9dThUKFMBp/zaXzuprmBCkEM1RMO
z/BaRspMLSSw5yD3d82F2FNA1BIdp5679fxpmPcl3Se+ZutbGmKe+lkM8n7S0g/8T2FJlAfEk4+r
T0GkBLMThqJBIBMjErZeo5vQmPYGF1DAIAiUTE9XzpBdYwZpsvv237N6BWeic6C7ZSwml7QnSg//
dJPJl/XwdF3ASdwN94WKDR+MT3MTv4XVTEv4ArcagE72qtDwOkqrKOczXrFGmIdtOa8KJt3w/J02
gYQRNZLm1j9zoMsR51Jryilfq6fdu1uIQQypeRFWmodNgMODbBl64LbMSYgVVKf5ZTKmZomraJ/a
iMufEkNR+FEXDBJVy9iqZkh0VHTUdTnl+jHT2RsyaqIdIfGOOTR63m4Nz5ZYw1q8xH0h9nvIFUdh
7ar8TmARgS+naeOpY9e14KLo1t2G9aqvRhJ0g3Dp9Q4BSYwDmJloc3jTDmlCJJC9MjXywY489uE1
6p+x90VRnahlRnda7yrcnK5/6z2X0H5bmyqXqiqAPFANEzigeMQLF07aLWuUEC8wqpZkTXWZ4gu4
i7L/SNzCA7t9nR5tRqtQeIZ0l6PDVL7YF6qEEw/DAidiun99tu9w5v6k8dzSzjsBqHCCFoec0g7m
IgrjBECQLmwUD4Q3eFj0kkOKJXWw8cla2d66J0QbDKVNpSZ9VK9woW/5OIYnZxVqKssoyZFd8MBt
sL4Ra9xO2u/bxQz8NtdSzv+EXp7YiyeeKvyyhcvLg2ypp3GHSNudT8Ju8V2jPkCOmZGfw+dhN+ny
Jc86bVhF6gIPQKwVuNx5vUxHbr2i2unXJg4B9FUF7Ol7+N3ttZuVrAHHYt4Tm0WNqyZmBbPV9dJ1
Yne/oPnEMNhUXuUcEuyjl5TyYgZjldFGHMbrK/dRFcZWy7cIW22J2bFvXV2xOSz6+XOFpiMAGVo2
ujovTn+Yltc5k4NhO7vpQk50DyL0kzemlcpz7HbLDu79Hd6lvvbruFMGaGZHx1dbbrwCB0vDdkaM
XRDXnWorVyVfPLSU0wps9mTD2n+XTyVBFpI+R9TPUaog9BdNj+WVQsORomkpLclH4ZCFP7my8DQ4
DSXkIHietv9+kqkyoUo630zPQ6nadxH4M0V2crlxidxxQGgzkqhVsdMCsndtdykoElGLdaXBJVZ2
ywTMjJkSp+xz8LBkSBluB6ZLE42W831VEMfZJEiChNgQ9vsGegwBz+EjVoiF19zbAH1vkimofssZ
8NN+Z8TDWdNi4olTV3P8erRl9g0UrrnwhUu5Fsi49FEXlYaDJx5Ztejc4bCs6YRf9IytK2wzcaXO
dnablw4G07lWutc0qDSiN+MT+AQoWXqOH1H8et0KfBVLZhG4peJdNMjyGXnfwimvqmCb8rp+EQiR
0p5DAHNoUXeZbK14YRYUOHwyBP7woEpfFnfdjN920YAsPlcRCqJFE47QmdU13J9fkE1NHBFHjj8h
SlVhMyHjXBfFZQB6xAo+Qurf1jwY5tKlzTM+5950+1K3wsqabeCLN7gv8IJz315SG7GiM8hLFA4t
YRwJYaY4+Z34B/r3gZiDV2WYzmxtWyPyRKZpAGmXh+BRu+p/q4lERYR1kX+WL460zbpbyTTxQ23s
KjAgexDxwMzwlzcyKNZyOBIthe6UM3kUthD0dYoxkpktwOI/KLONAcrC0gnjb166PxpDRfuhvKdU
ojD/pfx6MsNPnP9rHN6hIv32ZqmaP0J7/wUkgQXlXZbHmAnsiEcAdNUZ8bf24ks2HKb5lghF0iNp
YXFu2OmOV/4R+k/5RNw0Wwq5UUjb7V42qqiffepITGwxEu1Yt0NB68YIvpgsuUhhx/UqDCbl9qGC
qBv3WaW1pxD+n+Jmcs3X2sPd5CPq8aPlxylSI1JxUUTurTqRUlb/35RPqyTgjYy9xbmxx3OEtFIf
W7VQZKVGoZGo6bGUn0MqCObf1WhmEUFdObyK4DP4hswrQAsWFoFIVId+7JRJfMGqnTB7TUURCs+n
yB4dUoNj4ngyWeqOn8lanQ2i+swZjp7TDJAev5DaVIcnWwU/lVmt3NAx4syjPu5s5pJn2sCKGGKG
VmJyMMb4dlLFIIuheeuo8v2/594x5QV0kN19983dhYM/uy6U2EHB1tdOMQLSyg4oLvqFkZkXys+8
CUesGjDmmFO4748Hr7ifFzP5WRtPfbSELTmSU1lWcwroejTCCa8P9i5KwWhfvjxEXM0ePG9pVheK
y0fFKshlwS5srlzEjvmgkc9LFHszUXwzdSjGPIDpejgUdxYBJBn5hrSogquhMEphXHuNJw8n+ZD3
2qgYciI9QsMH/rIu8+RWSY83l8azIi+4iuptO0/TlXNj3ceh5jm6FXnE28D5XOMwwUzgNYR9FRHD
ggULWguiS8TXkrlWGaOfMoarR+ul1QHtX3rYGxkb1BcBDxnPHR4+44ThkdcX9e6O8SiX4IMDOWoG
cyQhKC8pqmVzgfSG3TWz2pWPS6S6TgBXb5NJBHCBvVZFey+qtMKu3y/WuPwSU3mD23WBOBo8O7Aw
OTq8j0a3z2DEsIn5FZSi0HD32WY81PzmY06U1ynlYUcl6xM7GkQ52/CTK/hYvQWCThTWSCWu161j
RdrISfXJXKpZae/z0GoKdcJguXeJJ1RtKPmqJoznqD8eCKzSVRhOmsNRbyiryulnsYJdnnSRNHEl
m1IntKJXS4HnDVZq+Wq6ibjUQEbBz5A2ZyeeO2BM6YCWCHEW97do9NDkm2oKBA+jPFBB/MneOSig
lhROJu12vK4orRxMYsb0T1Svi1ILMUlalHSOJI6jNA0AvHzo176DyL1hBdKJ81mmWvFBdoP0D7FS
e0lLiuuVbdwvi6mOM4l26VFD9FAndvVw6jNZSXQfMIJtB9csOyJYs+3aeZx9QYyNInKIWvVO5RZt
MrJnNGgIxPnVcTxAST7awl5a77EI9N5ENaAUUf05M1wvLoBI/xzyTvq2LNw+PciQIYZOQamoSk5i
8UIHlw3WIWDpQXtkd39fzo0wvMUB+xZhAiT2cJGs5hC+jULJi1mHec/4uwmf6M6RrXCVsTSP0VX8
F0SMvZiHFkhO7c7pyIcBZKbJVBmyoe0wLE3sxXDYTFPBXM2uEMK6yOA00oS7lHI2a8rIMtngR80l
9lJHv7YnUGS4q/zEbHH10Mr4KRYb2dV7/sx0XaAJ37glytuYyZ345PWUDbHLQ4r1tM7gp/XSIMut
PybwQ72VW5ctzAyHaZuzbV07bP/VL7AnlOfJdsr3Nt4Qmanjf3s4wnjX2YekAjx4n1cS7lMSfUME
6FqSWhlUzm0nM/RQSAyXrirAgOslcBvaFMiZEubp3FDZ/PR1738Qzw2kKOgRqutnprxGs1OV8h26
AUnJ/Ki70zhQTvAVfInmZ1Did8mJ8iuZsvt60A9UAjNtEW6FW8+oPamcNoULXxBV8QWAbgc8F0zI
2mE6ExvzAavyp7AmfcdSCoiKprtrJLebteYQZkR6r0RKoIZ044L64EpK1AGIELCZGpL8k4qO9P4r
FrZsE5gbJ9JTr1RNQOzW6AuIEJ6P0loAXaFPSaBeixCDadAqxuo+zol35X/vlGoquAlDllm02+HD
QRX2HEtrlyvcIMosXDl533j9R65jCsJ5KhBWfsfjelmG+2vPRhGZtGOYBpE36lzoQfZ+GZ908VN9
w6qT880/5djkVrAZDJdsyhuFUh8/x2wWvg7bzfejtYfxtLN3iXdpoBDG0yzayGsmlp8dm/I8nNPk
1X12FreDu7EsarFwC5ufs7a2jz3ZykIUaOpYmobvZoq4svfyMABSYla20laUd2/9z46E5XZi0oYZ
Lo1ZpKxaVM2BgH+67UwLCFu3iPykNWYToKNZzTRjYUd1wO+65oeDNDza1LL8Kg2+dqNDkL9Qlest
9tHxzgIV5m7VBX3dfmRqA7QEu220M4OFRqCX5PggtbUBSrPBIgzF2PvRg5/hrC+Nk9oflgicjT06
9c1InHJyd78Ip7UjjdctLR+a04a95GzVEpVNV1bn7UESYjHKrGHhDVzP4pzLeokEqahTJsisbgiy
j1uvLUY5p+aSUQzbtn3IOeDFXAFdCsXFdpunxX2yV9tCl9LsDEcd2+bv1tycI84zxg6nj2+A4VeM
YHrPJWX73Fo6swSWUjTZZT+QqsPd+pfhJh8EkTJ0Y1zPpqHGtDBBpt/LugHiWJxHNEMYh/oJ3RNI
82gRk1eS+7juyJHbFgHGCb3OLhFV63brSdw7jMg2VGnYx2KcUSU4GkSBuUoRG8tw62wZaBtJ3oIt
XCwvH1/n6hb3JSuvIFNRgbGh2PfQqUAoKLBsJjwtdm7UNFtuisCGS/TcaHJdKo9LvhprxNNzoMNG
M6UY/Vi7X4/gFV4ntVWyJ3lbh1ZzutaJLMKtCoQpR46i2o4uVzWWgGn4UL4xwyjDxCluQFbv7Niy
pwWVZTpgx1RTQvNE0b513xDx1jA/VO740pbVfiey/VKRAjeax7jU9qlpsw8kSPD0nzqITQJTkdiL
Fg7FjX569jsgWdIphafEjEPqC3D57nbWnczWEWbHAqiJgpmMQTelx+7/Dt5P8xN2Br7Zzk9k4hiV
a2jWCbgf8JhUgDftfSYDAhKNq972lQiRjEeELTOXaUmjEYSu44ADMb8ncF3PnjNDdPfvEDwTN6V5
aY45eg3gccX78A7Nh0HI+ccPXBYLEudENEYeQ1izn57APHB2HrYAHrJAu0NBA0xvgKrD/NIQTl80
Ak/mOLQGCUyFwJMMBRvjyC9INSBkd3Z1L/16WvZK2+414TMfcTbj+qe9RlAfi8FJuSpnOjhoYYJz
ZfH9Kc0C8YaDgVoDGMTuH7f4CCXDL2k0CZCeMDmlW9IfgcSdx5zFbcc1dIKgnknBEglfKRMEpAz1
Ei193uccVSN23tcCxc8oJd8Jj2wRAxa3xA2/nWWAfwdKpjVJbYn2w2X/pBcdAmi1fOCWzumtS/zH
FJN1KeoNlDzAXMRwgqptqx/KCWfodswavOSdPQBXP5vgHleCo2xAqwOm9zU1+YW1nDN88lfZt9k+
U9kCV1un3ulrBno184gHRfdpkzl0WrEQ5Hzi2ngIuXlOm8cntbF9nPIRo9L77GmBVZ10UyhalMOW
SW4nTKX5+p1b0vebR4gVaOIuUyBjsMkfQMUeI+EQR7lksiGb66NS8Q2YlFVNk8f0dsWXKiY+Il0e
Hqz8fFeYCHEZ0YlT41sjwat53AhHlCTmvnFhHRe58hISCOxb5PyO9BrEKYWALTIzF8UttBrIGWjj
VKCNXYShMRjvKoyfBQpka2DCDB2jtQDzPfNrctznHra4/vII2fOfdCrp6oM/NZwtqoZZU3nMMVfI
DtqxiYksB6H8WUMetZNwbRctGrAq/RCgd2HIPOYMyx5xk0k0GGbVW3JaQQ0ZkEBTKvQGupCdLDK/
L5PsQN7q5p9vKh0Ji2B/Hx8eehuMIkaPsxQalin2256E+a57Rdrx/cCbisAQ9H20GUP6EnlQQ9Ft
qXigT0+mki58NxeBtV3dFM9o3Rmn8pjBELMDzh/cINda4Qd0kCp1KBvWR2aU05Dow2udC/kXDNci
jtrQbkQutr5Txy5OxVH1g5myZfduzG0nWn5ALk+/vUpGk0eFtyF8dlh2wVjtekhZG/cfwL3jCLbw
0hg5boQLDDyYcF5m+rAu0740YKuDyAH/7j2Ymo7QG5qMqqQRXkKfYO1fyBvFUj2jqqiqu/YLoawx
Tq+y0e3FhE4amKUbosbzZ2uhyJ3fAvHdSkEitYegDax4GAk3oWIfUeuKRF+RDia/P8xrK7wroaiu
x80rTg9z8i2lF+wTxha6RwgGLp52qEZ7yyuHyLbuA5M08dzEzArPsylBMoAkOyn5O6HiBSwAbHZF
DFNkCkRKQzWpM066u4FnddfY/CnO5HzMKFrm/0kgwFZx0a5+Euc5FX3vQ8P431ZPp+g39WK/YQN5
6uDeZzhunUFISD5tSDhp1ozekMtb6eg/wlnSJHfMTgUi0ixE7Ffum4myJLieRn8bQDcYqp5ZBOl7
hPivFKCOr84E2aJhhn3WsSqd4f1eQ8Uke9RM+wxpPcV52+pzBa50upJs2+F9pTv5P2lhkwQrqOM3
AJEhMawGHbc9Lnu1KDJNtvy8d5uprPxbmT0LrH28duLTPiEQXJpTpS14fv9j3S9u5OX8TEsF7OxY
N13QQcESM3R5E1/pAWkrn9VcBX9BFBB7B2VqahR+22FrDmZr/APs5OrGnE3ddzvQvhot85HKoYjG
Kw9y1f0nKB4JTkVuM0g8bRc3GJ9S704UoyZ1RkkUtXYJtUyN6LPAn2KGiRkKkBSmfEzZPS1X4e/3
5hR7upzBEzfHAasuzWz15fOVdUR+1cPdTMvUo5i60pwJ0jI29S0MaW/u8Y9O9HAreLjQ9Gn6utzM
TVaNHzxWeYPlCGBqVET+/HGSVEas2/2N/ttag/AJuEpyfEQCqj2X2gwqvUArR2dKW5JfvlZxJ9E1
6gJuujFkeU87J8g+XSRizdKv8Nk54RaoKLPhAOr1atAy//KVvnq0ct6hMnw9j9udNyou1RmB+o58
7kW6i8Kk2hnu0RZgnUXP2lS29ayncBn3Z9VpSKAsa08mynEeUXu60TUXbsUViSTtXxWEiJfPqT0Y
dctlO/XJROw359Q6HlTkFoCOkvZtdjR+Z1txkMeDKYzZ209bgw11awO/Jkn9n8lfKK7UprZNKucQ
Dgp5c0ewJnukX2JE+vOGQfkbwLK5EOn8Mpc0+KexiqhJwATBHwezCmiuVo5aongmZGhNYfQCxZjm
+w94N+4hrVv5QL4VsHblRFEAoUXmsGLJRxljfi6S/D+vxCjU+pFLfLSgj2Lrq9QdSfCqxm4vpiOW
aazDN4aA6r1yXG0N/oc8MVLhTmUzLx2NyNSzaQb6afCGs6rsvo8dfFXI2Fjf1EGQouixPQVQmbkw
RNtOiWCV6GN5Fz7/kZYqbFn3uIlmf/TPkD/o+Qs5wW6YQzJUe3HXrnu08W5K1+FXQJxR6OBKvKvp
N7ERRC3wxG/55iDiTRGILt4vkLuSA8ZuOC+BJizHHE2W42G9kYqzqJPkQvM5s0O9ISHKfFFkH5Pq
eBTSBjKZG19Inwom5EhOPAVP19lgwh1mIuZW5iAQ0ycevkycYYsSOnscbWUA6ec+jF5tYpFMKw7n
tAUjAotGYcoFw0YBKyQ2XJ+rS35gZ89x+ncRl4j9Nb8m6jsOVw7B/NtKQrl3HOz+6R52sH74v1ro
P1kH1hhw5SsXkG1w1++9MTQdCtf3VvlFfynkLjlG4FhAKYYVRmNtGeoB+srU8DyIlyF0oS/tkoQR
/2WawD8R/lp9gawWq1BYM+h46FrK2UsUVi0LxoxRuL7AOcHJn9nRta6tlk5Z6c3DmFXRl/2uX5pU
/gWSKauCW16xN9TVoeZlCVQjKMCSZ92AnWYnBuY37vjNHW09Yl9pmi1wY//Km/G2Ntiu+zxuTTmb
vmY3TfudDtjbmkGsygsln07NVQI8TfmmIze5tS/0BXTPEJIXFcA0/5tGnckwMq8dpt5/vL8oBgLI
yKH4Du9tBt6rejuSQSI17N0eYya73O0hlanE5o2Whl7+Af3Qh1AglhZaqiWwzDt7pAZSmI8DahwG
HPAtt0uhAPVmFNiPU+jraZiMg+2FUGxfwFCf3zfQ3elUXYJnO92hq7GaM7kv1rNj02Dje9x5FPmr
WgZqpvc5Pp8/b8Z6qbfeUrQ8Wl8TPwj975HYSqS0wEo08xw1OCir4XlwzjB2ZpIVvoh2URJSzTOw
yjbEvMFIP8+ek5mxHVw/OG2Vv7iFr5SXsy7aSuVn6TfnHlZsQ7oaWh+brEOLnnBELahJcBxRdyOw
/nEOyGwQjjbT2bvkXh7CMXfhAn5Gc7foGl2zSzHwpf168W+TWlfAxgvy5nk67u8/o4RrQheQpxQP
rVKLNlUDBUQefR/MVgqtlJXI3Z14QVU+tPjy10sDFKkkS5OHVQSSiFqVQsrF79yuBcZcBQOZyoAD
xQu9kf7eCUIzsIHJEUOTa+9wzz9PrPlj3gctobgAoPNxHgDMblhQ8qnkkroCOczMG+UqaBEaPw2C
B/cYbCUzhPqPsiLbQneUtUtPPTQMbuCcqIdAboA1jOoAG4VW9I0yCZ4LCrTiXyhsJ3ZUGybGUmaC
a4Gy91H+y9PQQk2JE9Hdno1II5QH2QePNuGkBJf+O0CzFsWjhjpeUZ8kmMN2J3ppHqJ8LCcBIWBn
yxaA7V6MT+ttEGSapvQM4bT6AZV+szLHrNjNC3KvUUrXPrX9NEh3UmSjPKFy29goNo9Q1/5ak1/R
NyDX7DogLWNHwYOt1LvtccJT8DEKIhy4uzNW6nistXHIpEkbz+hFgeOx6zmeRVHelbH3gE0F49eK
Vxs7elH82/Rr+gcaQSRpuKLR+lzSFtfgdHoslcywivYjCax+oHVeqpO9luS4ior2pBvvwrPtMwQD
dXLGcscMWjR+i3hGLSl6FbUZgHe2YMgZTV3ytWyqk7a3VeTUARbGf71I49nltUKdQsSmazVzpKjT
JTLLMD8atGEsC4e2n626QDzeBZoDc3YM6XRRQc3NxZHlPUwPLtrcRmiL8C39Jw9XrTdq9OyqFbVs
XP3DXv0yRbXptE27ZLmwvEkEEWgqdL9i25rEnKKiI2CXFADmHJ2hUwhMsISn+u+23lBchnM3blil
sOkMY0VTKnQIeQh9ZOSpJkWX25if0454uiLIAelHyWpq3yOc5EVk7TNHqY3i8/DeWu3XU8O23ghp
+1YcZJMQKcWz7/6qactvXJISO/HIocRwaQ3EBB02zVHvT3rGjMUiE7aEEQSFCeBMnFKla4l8a5rf
Bci+NUv1dVZ1Kj2q1EyDespRwPtfsMp02NtXnZ4dEm/dI5QkrlVTqhgKAMj51ewx0Bp34CF+U+td
DFhD6a8g0nn5gG69MVZbHc2htmxykcYa2co18T8IhZT1pV1eA7q2+gq+HzL/K8NyaJIv/5BELK85
pWiQRa8M04lg3+F/Vdqa9rbmrJbSUVT6n/ZEE0u7kHeLl9x8Gr4iEC1pmCI3DezLxRKYNZvAMh7f
QpIITwG+oXkBDkGvj5n9ryRAwPPeqknY/L5VnRWMTJC0N0toRbNI3N8Bb7mvqgjmkLKif1BFDCpg
PDrCktFxb7UOShh+fKsKz8rE8P9sk7NPWVSZQ+Bqk/GOv7E6n7/MKbrAew+gSsTMmo48RxZ3qv1B
6AB7SDN2j9hMkq9qQUEqn40OaImKojRgImQW6LABl4kw6vHpTuDiLYUhKDbXmrVdmCSb7GxcsHrF
sreDOOrle1a7vpU7duboOfjY/SUBdCKM/W9tH5YkqhDiOJPxc6xjdvZRBtCpTYSQLC+do/BRhYXN
CP1RNkbjo1OOF3cQFoIdRS8kPsriY1tiT7y/Etxmqv+n+2UjdykWEjigdA0CWeb1Hyuw+zypZshH
bg61dAuf7KAOF9OkXx6s1rGrDgr3BHTiGuRfl5BN/akjbf/mPvchDwadWyXkvFNha7WT0hUKNzdd
yC97dm/9/pK+wV59kAwdqQmFjdw2VCIxBerfwzikB9V8Tf+VExfAWU3iQDGdsd898ZrKLBC7yg1J
xd/8oWNBP2ULbvMR+KU4XCgntUXpNSFZbCm+iI0MX4RLWAYNBwdJF3owyTy2YVMEFDvSRBnyIPfR
h9kcCMZxw9gLW+HPMOCpDVbUsN89iWAnQN9i5QlNVECZAFwXW+wwq4ErzgHlQDg04oDLVlVxuWx5
55SPLILvXs9QIwOf33/MhUYJn7R29s1l6y7IzDuLntfhCXgoUs6ctLBqEU/hfPAJtrGgPNbEX2em
z01EOv6XmPnMgq2K5gEvbd7kUjtqTsCoWl07BnTnD7PsFxYuO54iaxEuhG6JId2dcuVpyzbdFeuo
wPBDatbzifgzdwSpoxJsa0Dj8dahJ+cDr/K/7sPi1z3D3iOdYyJdkW6SEuiQASY48/TJmXgh8YUm
sZZbC9vpEZErNE3i1Z15rJgidPZ1R9Y5lvKj6feNCPjohTEef1g0/q4KXcn7fc7+gIiymoXFqMxm
+f3k2oaYb+UkY3eRlzX/EpR4c1Wm1IeC/IoKR8ELR41ArLx18xU01se09PwbyJGuoXI2wNt8Ha/A
B/LgG2yqLp2jNISxXbA0LhQG0Zry8Nmrw1a7d5VMVOSTvAbhSXN9nRHqjU5nAGG6h/Zr2UbOZRAv
GNnZ+GwCFHJ2Zp+xhA/ruRZh5veX0NMNBIwVYfojtPuoVFIBrnad24je+yNJdu8/5au8RYH6XUlt
fakKkhoYWPbt5BbIz2yS53pA39sXbYnh/VRUdGOC/p5M9BUd/4zdXlY3WkJh2lu/4C+o5L2Syp26
obEDoSy/ILugIJKNKPfambw/ly6bpvlzbEKC+VRY0SIA3z6WGtSKuSVQdNcfnouNqYgsbTwwAq6v
xZef6E/AU1p/CPYKWFmT90PoB7TRoTbgWemYCJ+ZyZFpsJs4bz3/mj1IoXUQ695ohC2jGu/OxRhk
Bsh6yFfozQOqknw+gFTgNvH21abB4HkoY3UQm60kW2VmbaSfWaMbJwOUQmTrSi0m61yDIK1Oh7du
PA342jkFKPFB9/WbPLpPo5UbRp7y0bda9Dsl//F2EBw0HNkzG376b4FWaxYPVvT43Ixr3arwDVvc
Pq7dZbAYUmGDxGG4JSPLlux0P71Y2bBt2drZ4E3Oe7kKryku4igqzto6jju+oXGqnhiVsVaa4Eqf
w6wfd5G9G9ye0Zh7Af74x8dxZB0qOfGnQa9LuKF/scj8QqBNsSZgme0vKALilUiCTvljRlB1OKYF
Z8VK8CMnQvdYZnr6VH/S6efvgPSOGrCSNAWf94s8+KugwrEwfb3czd2jizv+0j9UeX/npNJ9c7Hf
WWgGABuXTKr6NnW/elXhWB+JvN4hjk5dvt/eceeYC3Xp34w36jMOQN54HYCAyc+dGWouCGUaRosY
xc9Pjje/vbYyyVU9VRIHBunRrX7APBChPKCSQ1j+gWEBGWOHtZb9K2nUrrqek+YOcr9f1/N9wHyi
JUyHzVZcNHG05YZEgj7qisKy705RJgUxqPFDgVWwcj3KLtIwP6/D/bpwItjVUBrFtVL2sYZ0WtCn
0cJC51x+eQy/uS6RPpkqaKdfjg7bxZpJ8mdF5EaOFHc+Ts8oVnv0i/sj3K2t1tKTNHZjuWI8NBu0
wTfitHH/UNwsws/nYt0pYT4lT8sx8faI95psjermKEAls5krx6AuieqDQX2ZV73ezC3N63HWtwwy
Y4yLq0y5wX4ejT6ftCj3T/IjReLITKhMqER+kfm3MF/XwrunavTm4kkcsXisbsvksyoFRY3r+RK2
mfV57IvBFj6N9SgJmpM9DPfm1F6MSDoQgq0GFpnOXDCh+YWrfe3M2jXgA/UENCeHvKqxQpLV1x3v
+vl3gcDLIUW6XlQ4C80e8tgvAWGhMIJYWTlLV4o1MvTalNURcj4Vvta4sRE/pvVu9SV4d7wfFcCS
P7OjF/AfvCQC+8QOfh7aR/e6rjnmuo2eqaZLKqW9rmUh32KN1rNs4dVCqDRJoUrp4yUOOyKMbiPd
Gxilrx+3oU/dHOPch/kxuUTudb2uQIvtCqvJJHpkzJUPyfMw2eMHNAps51UVdBq+3xMlWtcDLyOu
7SPzEisIXjqfQL0KRuJ150cn+VBeUZ4OkHjWrl+q8xRp6gsteVFnYAQ9zsHWTXIOyUIZqQdGYZg7
6e0LjkbjJMemNkRp7hOXpcSqHFdjps5AeglvKpKi7FPRCd7lvehcNLJMul/l/oZsU1Fw5kZvjoqo
qxFONavFqqfpy5+sW+T/GmkjoFmlUzjsV9FPuq0B+Tlea4rgLJPO/jtnHrIKFYyJhePhepkNfW1y
JWHiKIL7ljf7IXAJvQSYMOJwOjSmDPzprCfozjgj9sJy1Luy/1vANnZDJP85yZ4YWYynQQVGJrMN
PZ4J2EaWfIrMLwVtRSBhLajmnkfZML2TTHJLhFYN+sbkZQNlkE/MXf3Yl7kTRV07xlRc8hRroqW2
dYaLJOtOlWz9YNEDzwUnWSKNJ+YmZzzG1AfNfjScRQmpdZZud344poRjfRkst6ZXFYwwuXIljvhO
3tTrKQgnVs3lSOuRMI2fgWqxCGCYO7AbSg1bTYnUyCbWx3SYjLKKzZ68nH0K28725ihy6ar3lbGy
eKr/LsTeEE1bFXs/T4QfxaMgyUXrSM360svLRc8Gjy14ejbvr8cYAmjVyuNTWzW5vC+nsLhrv3bC
0dSYqLfNgVBnxmTNvPrhPVKEIixVwiqM7JFnyxNYVVF+Bc4SaEbUEn/wfQZUA1qkAjqyPL+Yh9zE
6NXoOzLx+5r6AL4KOjxFGj3LdTcKSgxx5B0U9sOwPepDAaPFw65sSka+eOKDCXTvQGg2SINpiZfj
o66aey2wXhERnF0tXrqxbMBWvhO2bwBycplF4nKvvy6RCrI0eEgHymNQnpH9zQ4y6jbhdtlJAUzm
Mlkf86aDhJVXvP0u/HnRCuomA6NkgSHi3fz7gW84/Ea5Uy4xwArB9440jj6Pi+WlxSGuyTgoHoH/
exda2//rNOmvTpuuh7zYO6PbD+CWA/MPq0/hZP1LgHsfpAviVsT+oTqeD6a+zgELAvhKkhV/1EcT
y/ch7H82h5EHqItPtqrUx95Q7GzgHXt5NyHD7nDDRo8pbB7wrQXB0ugqv6/96XcywXU9PxPZ9ACh
1ZqzRniUkfOd3q2dGiiRjAHghatUouVtdX/JFU+glBbqSpC2C5p0cDIEggGjx9+GJ9AacQU2PTKM
wWYLpYT9D8Kxzg++DSX/CmIbPlqtb1yXddgqsDQZvoLJqZOp0oxlQZEwFfP0DXflQaevJwaIv6mi
skOMw9JKu/MIU1UOlVrK+D7dPPWPmq1yMyKVv13bxqlUwSB0iexqv1/d4BcYJatsKoyp5PsGZZHK
Z3LGW3EXiPJ3jVYkb2L4UZP66GqPxsMPG4oOGdv11rYpE4tuny9qUu4xEa+iZ/7CRSsXssYRl8yI
LfE/pE37J/9idxD5J0yFasue0kFvMW66ITMkxNKHEDHENyYbkykxJDxUqkTb5+TOTUL4TVIlBQhQ
r7wo/BegxHOzqf/ojnO2E5yb5j+kdc57+9FVgpmjr02SbvviqqIsuuFPyxq6g3KoKwj3F+rwzAjo
s4FyNUDeGjP3j5xCqrSBV/Dhci/c85YB7gZkVKKp8+K8576t4NinwWJtAIGGXCLGLFlu07GoxDBR
yAnwyKKLJyZeU9etC9ODMy9EjycPCjfhJLSzNVNRhTLSu/HsK34S3PRyhxtGOCMoLXIb88/PW3wH
MnG2UwKc8WrtbRO6JULMk1i2RaAGWLNTck48WqfQLp5VtQI32ajzTrH/2gWAYjHc4tWaik13uwio
2m0juWZAdDUFqBGzHAmMbeG4XeYljRg63EInx1qH961lEa3y9hsH5zGiIqhaQcEKFqTWKllKXSNp
1xUfKMmB75JuywyGXUDSEuUc4djESiraCNJmCtBD/NICLIgumyPdE9q4JOXqxmDz+RC6bP2spHZ/
1Omf7ttYlxy3dGo/A5noxcSaDcnJYwsDxF8mnYyvpAqj1m6AXVwOcTpSMLGFP5AR4xXCHXVftmbw
3UttwXfGall2UfH21K1cCXBoQcoU+LtCfVXQ72JH5P5WBraJCwkbrxAXF39LzTW8en6X97Rmce10
kn53Ctx/1zn/g9bp5E7XKTIYKpwjX82nm1h5/gdMlsSohtAE5weUoE7E1f0rDjd/kkbe9uZfH4xp
X2trdfLBCpPpG0woRBZhl7i/BBsw0AqdLzuX2fP8Sdpl+td36cbFaAgpAMYdu9iifN98U8CmR6Fd
1HMlXJJ7O5nJj6Z4wlHotfcj4Yz+BVAV1IwhpktkyvG8kAxn3OajNArP4+1iAjvnXxh8JEGHoeax
4H1CB4CvyjxAbUzsUzvbMFHemQALpE8YhATmtNb0U2ow9SXXJwmqXcmE1UqO++amfSME5o12kpwk
kjoMbq3BN1CzPv37QO64qRvqHGfnKdN9XROds3ZuoapfgTAsdDTzNeZU6CdVW/PY/yliYZfagP99
OU7eAk5AUVyS1IHgWZjxm/vU5ojaVk3eNDW+B4k01iK7D5nthJ01jrjEuyS2jNwsV+1ZYqeOwmtk
0MoUQLjOj+bEVHk2lWcB8UclLIkBZb4z7xAz8zZHJZ2EIl9ZMa/IJk87pLrp6iiqfQU4b9SLV0HU
tQ8PLbHsWzJmJAOFdRvXlaOqLfQZH+52mid5ZPMD/rmrfC9fj0XUsYbGmml8PFLnevmag6ySn6Bd
gm40L4BDRaZB7G0xu42ry2hAGGZ9DZanx/3p26kWbJQA62H9Y9WwahWecbR2AOKUZepJVU3drI5q
KWTDuQ1r/XJU/4L6wu6imEVTr/L7YhA5INILN+rdqYxU5Qk9qvKd4Dq+6cTkMAd/PTSeliHL2Poq
JduUjsxV+m4EY19pq14HFDrh+DCxGDHe76odTFpURM84vVgfa2wyxKhtr8MoJU6eFnLR21Pc6/nx
mSftFNMlHcstZt0AMMAW/epEadyP/k3OXsNMR1kzC3Bzn5grBzHT2glIzsqxzPsoT4FCARzHSyro
KhdavS9Pt7WcSp7U68yqaSNezWAE/kR7rf7oIkVdBr6ydjmcHeIelkAKsJhgIOHRtq/OhP1dwuAK
DGSE6YFkFK3dWtgmKIQ/NdS+kMSyCospE4PCpqvcp5EH2iGR29+w7uwI/T0rwsHBy6UtVwQeTV8G
w/ImvEZTpx4QasyMtXsnIkocRVbrfIxikHBdweGMXaR06/6HhYYaePBEJ3SJCg4vRkDsME+HnYil
mV2oCl8ufECSw1vog1F9elUOOdlsPfA6D619VqZnfMLw1MphIpFdaxNMMmxKuzHg6VFUqnhCL+gY
Qnj//KWiYexvB+cbxb87lmNlZp8AFw9qThRv1kZgfkEIGvTLTauhiE15p9FMgooYs80XGhx3BDuF
gxaQd+5uFGIYCEtGHN9iuEY6CkUuW3rFzhlnxORrypL+xnzHgX70Oc2Gfp5TmvSw7RZm61Lgc6Xu
SksK2u2pOynV1jJi5cxPPwTw3KsfHZ1RW5qTTF213Hf7FUrBBab+7Gc3EBEHNc3yX+iY2vL6bFTv
hTEiT12iBTMpCAVwbVPtLlRaaNStWXPwVvn+u7mPi2GSS5oBAvcdKHuKgsxqweGer+CwQazbB9Ro
9r6EnK2xOuIJ1IBUFdz3TxiMeIvsHUVvzO6Im2dKFHk6w9TC/6cShpdDZiP4/+368IjDAeUGjwMZ
b5kfbmoNP4xRRUyPmuP8/1hNuhgbVVh42fAloZnCRJI1gx0Bi4O7dsOZLsbXdhQsoE9cK3MMCyBJ
V3Emwm/QmITPTtXMGqCwvTm1RjCTcaPIlZiUgc4ey6SKOTLb3OErqNGrvH79X0m3Iax1wJjOEu7J
gofTsmHNx22VA051RTvGPX6ikvb6G93TFGRJeEX875nsVjGwC7PsQ1RGdeJzsVG+hNJPs3y2aJ/M
L7SwwvXYtliZljOB3dJIX6Zj7vXU1EYA2wxnCrGPaMWbE6upxTA6UG7ziHaN0RVhy76XpXmKU/jb
aL/H6FFOLxy1mlkyYZ9R3BoYbwVqv+H51a8QkZlVfNz7ULinf3/Xt84Rp91MMYCAIKLCmAt/5rop
tDtAwEzTNLWlRFNdc+feeyHQISH59HtTHO51qLEBAR68CxM6rAsmb0taHUFqO0e7Yv37Zm2NxZX7
wonbqfBgw4YubZQWdBjwpk2q5WLvYFFfpUbTMaJ6Lg24Zp0WZLo/rbBVlW7b6cgDdpV+SeRMYDmL
zaBa5kxPPBc4YPPED0DOYM+676jyNhE9G9FQyJPy1yLmZ3VMar7+URI+c7RZZFkA4KFLmixzHrf/
mIMkETzbSO2RCFC2BR4x3NmuPNQnQupoxc246oapL3IbWjNqeYEQhnS0CB5E4AaNYpTgdLULoJ2y
AMvEy6H8DiFlIeOAiT9J1pFD+mgIn1i2I+mwXgO1OtvcFeL0/4Ixtu/hAOgA/L7MMoL6i0rfqqhR
wEM3jYdYvM9s4rXHWstq2z0FtRDwNLIlISsfVa/JHKLwAIS5HQLaq6iObwQBGVHRT5x7u8m6Xr65
3/zKKphdEYSsyeYWLHBE6xNugsEiACPg8pOjVjQltAev69QjCFWzGUa/HN8k0isdbD+G9Pc6Jutj
GM9GiTpUalxFJ+eBo+TZvlHJFyrLzHHB7oDoPH/ADI4UfGO84j7uIwkKr5VVS4/sxZpNIZ1D0Qfx
KhAZLugXH/nIfbIf5CuFS05XF8G3nD0blowu9TqIWBzNbDzJtQP0HWLTwx+96RAosnJuBzhgk/hq
RmBENp3wC2vgJobrUAXnHZub+XJrRcqrvI4Zu7xthvoaHV3EqBGB5+k6X+CIf+Xwth+gpePXO9WH
Tf1T18uzX/SwCRE6TVjSs++rtMLpsvx+SmurTobmBlPhDXrVALJQ8pzpOvH+ojOo5MPcvJ6R43FM
KGpSCRPokiYLAntgvhN2kHX5y7m6krIg33ukSoShdEX5j0wpkfz8dMjWDypsPkTK01nKFzr8CaeN
q6grhtEitPBfnk5trlUe//LjpiR+g7NwOHOE9gYXfETbXNkFDzOsw2zInElC/Fcv7mSidIYNm0zC
AXSe5rtPi/mY7FmPIRjR4OSGoe5QMVuv0xFXLstAyOhTHaiHr7xvC9z/UNr/mANjDzj2Kv5p47RN
HhMDVOeRF86zg++Aj13nOmIxWKLSUFut6EGF3pXgFCsS8ZBeB4AKGqFaXZUOt3SzZd7uTuVtaII7
waWEluNCDBd+akFjIjrK3DFuOYNMOVCtnp0Zte3icK2ICJq3NGoDjT9k0CZjJ4K+cY/dBygzH/VQ
1sesdq3Av3J/LI5nCcqXwjojrD/XPRGZ7rlXAdudRR8Z7jbHO3d+flLjCHfc7BDQEi4OMO5xw0om
FoEJjINqlqpuu5RYuSnY53uytuwHexpXojv9aVRWLrDlECfTp7wbIdBBytI8o3cM7y3teEUdM884
npRjhB+VZtfgdR5fyg7aANeZ6bx6q0XaQ7DALSQyxS7l7O9MCKsdW9t8rV6HWYncoY4Cqv9PWvHb
2/yNKE+zQXrOhvDy5yyU9uSLuasFZJ4gaBT+KTTxAwBdG8z3j1YOL7salwLw4m0+6kcqC2prn+Lv
UPhrMPuugsgDcib3yOM2U6/3NaNIN1mkpvsoJ3Svch8ytrxJVBLPaTswEo73ud7lRSqTPCLroifc
fsHaovoqtchz9QkScRL4ikYslGWbYvzn74IK8sMwIkM4I6EbrqUd+6wDqwx93sC9uI2LVbm2xfZj
0ympb+y0Tbz1LHb75g8ePkzrXHND3fzS88gtdjCWDBpse3OrfO2QKe0/zYH+R/4NULxDyqTPzgpf
OCFrx2xEjCncNTMDgvIcrrdg3ICvkCcyNygGLp5x4PNRabq/2RHI4XKpyhzNUIEQoHLGp93mhmpP
dQK/KJHGriQLZuuIghbqyPS0lQ2oYc3CBDqxL+ek8GZI25WE1PehNPqf4W0gxxKEEkvPvfBPUbeE
4zLUDADoSbG0bm+S03UUVfoCZK58tIvIYRJJ05UqVc0QDwTvcJHag4QRml5i6WlKXe5VC8usqPDW
rFtDRDHM4PusxbTLhtZFbdSuZNxrGYA/ibGEYekZSKTXl+ylJAc923vqEWWN1qRfAyakBRFch/y6
R6vXmcKEu0KvEAAqu2FyzGBl9oKEQuCVk73V3y3b7b+f44FrNYUFsChe29ZWksTQb6NA+UYNcvG2
YL2uO+S1t96gneetn+gqA4Dfm+C7yPD1NRvKA6cIcSHsBIFnUqaK1XVf0prEvePFjDg8hxRw0r3V
YR5E0wwC707krg86OiMEdXpnZ4fOkQw6oXKP8NLCjkhdWiUnflQX66fE3+NJyOgOY9dK6C9S9ZK2
hNdRZaEQbBm8cJrimGkKwTccfw0wrD4ScTCrGGJJbpSJ7vsyN3e+ijSOdfrmOrY+4/ozq7Fg2yo8
KwhLYwyqB6VxAA3USUVbFTzgRkVC9GgqjGJR6F1DTcyHVbw7Kim+J995hm51yQcHqdziyUPKqTrS
e3x4qEJzbhkruF5odRmvDyRipto0HwrAVpQz9/ntkfGk86nL8bxnCApax2YQNojBVQ43uwZEsTm8
IE/c2U2Y8d7cFS3FQi04ahpZobW8l8n2EfdWoCJpL7xK84pQKbi+Ci+Aoph8FJc0nilZsJ8ouVEJ
LGWhfH4+HJo5gAkF4rutz9jmJ/izz7VjoKZO7MvGjkNftEYtM7N9++NWuq0wYsnfOKeSgLQ0Mo4I
M/FFc4oGU/ePsaIMCT4LDiEm6v7ty/teq2mxnndWkD4ORlQ6vU6rRfgN7rxs++sYESkUL8Jqzogi
1+DpHcjF441PIaFaHdqpu5HsUMyDtCGl5BZuaKLag+KaSaZxDIUyfP6BSNKNbRTiYQ5a1Dp3wXEI
tSmCQlcN4yj8JpPrwpINIP8zeiJ0W6wTuPfZd3ELhXDajyUTUmMovQRvmMLhlfTiBEXnBxV3ZiiZ
RGL4iaa9qC2hq7YmgP9d+Ie03qIOcRtZbts+3obCmEWw2yEob1iirXp3a5EM00UdGwigftE42n5r
+WocifnHs6vNO43QlPyohsJZtoMJ1K5NveGUABx9r5s8Tg1VSZUAjZGReOtaeLAXhx4ua9Cic3V3
S0Ee01FcxcZDPVSVXk3GElljEFJZ/lSxyX9Yn3x9p6E/W2WKhkXG8m1x7jFrQqOZRPj/pfNIluyC
Mq3MFdk3WSC5tt+0NqKF+JCr4HE+eNtXqjul9NFFC/2AL2VLIpVagYUXYMC36kVb+ZsuOe6IcwEA
ZBTew0q9NGDqlPwWlvRe+tZwi9sm5H6O8EfOU5BTsxP+1ruNlSL7vY9aWfIYq4c6D/2u6OEh6DOb
So8ysFvZHb729/2cCqTMcHdrCbYUHbllRETGgcnPy3Mxl5S7oqKa5yDVfOcI3DqpAWPVsC3HFBQ1
bYGMVelIB8Zc5lWLU+lYYF40pGQsEQjh8HqavOVBzQVKAgq257dPEC5iyPAHDH0kEo1TqQh0V4U4
j/5s1mccoZQ4Pu8DWrdvJoJsue3rO1NIzbjkPqjX7nUXqEWBKY2Oktk39ZMFcsMuhOznMf2U++Ho
29UWhlXjrI763o1nF42DLWi5gM59OjLLdOERDKmz7JsUcTbciPw8Ip41lf+nWsMP9yW8X2+DE21b
s/eHfzbhUHMTxcCwx0vxP5erjCoYFfg7jWSpV8KKfdgGJ/EBG37ijEI4D6gEuFHGboCVBnzRVG6d
p6DXrhYHUz7+mmAaB3EWr/x6Z9E7+s0klW4v/ZTNfXm1NiEmqXXQUJCArQ6WVh/VQbe8o55O5JfJ
B9gMtd77CiDhiqJR98esrQ8Nce/EkFhmQCdj9zQuWYBPzVS3smt0iPhGfpJAbWLwUv505Xyt23Q3
BsYJdjT3gI/ienbC7PxyWPjl35XijEK62jxuNDuAtX/aLcO6vH13LDy2AG+nUuKgNpa//jj7rtK2
XA2+9kvu48gRkhvENZxL0anZr28zhNjcmz+xaPwEIupGD/1lLBbfdfKpKiuZ6ySD2TWmBDDMet/6
OBgyHqGNC749pbuA+LOFPsNspVndQLXRLXvaP4zssW8crOIZRMeSv98axmUhDyFa5ecybnOY5Rhr
/ScxEsJnFoMy3OVEri568wzC7HgcP/R8sGm+yVbHUTquagjd71gAIjQnBGrDTaQgTC7Pg/dsIMPC
mHiSubEeEwrZ23cyx32Zp04hZqGCU1pqN3rPVFY+IbjJAdeojIrjD5VpOawRvNG7O8XDtXcUQb+H
R+AAD7BPM6lrw+EUW5CFpjO1mgz0bSQIR0cXlkmQGwCEJZiZHMUVgriaDr88vd0VObol/A6srkwT
/59VuWhEfFadmB0XgB0rDxf5ENY46RBantpro19SfU7QEPeQmw7UI+6bP5Luo+vgueQoyrxiJR3C
Q07PSLC8GhoO+d3PbsbMHI+HU1rnaQlmRPRvYUe0Ck6cMWJo7WG/sm6Yoey+Yr1V8F/uCh3Qmfuf
EEw4h9zSzMg2NbDNjAXey6MBZltic4EWqdCfzj13my8gzY4flCEHtYJmJ3He3S7CHkv5fuxKilNc
An70RRRm04u4lQkPMvusvLTc4ZTpMxDTxE29hYLM3QS6leEDLo74of8NVwxbrObsVl7OEMpin3JW
fQnqjCbq++olPh1Ry9S6FxJcT6g9Q/YcP1eLNgtmPyMvFAOxqE6mjBmAfHJlo87XHadoB2RuKZKx
ySNNHtBRpXA7CM+6fZba5lGlBpN6jHgQpKjijOYvPU/PZ+vLbKsKIh8yvUR5HLTQShKd4O5NRRQU
3QKVPyQtuH7LWfKkHlm2pEgQcwXXyA7o18mYX6co1ddxheGgGcSQeXbvesaYGEHjui6NoAt2r5KC
7Ev4vU2EbIQvudBWoH+QXM23HWr6Fj9Rcc/Ha2bpc+TWQoJncyj1LuTPd6PpECajeQWOEIG46beU
vLKrHP/UApKwpRwV5QPZsRs8zLdJ9kM45S0WARE/tvkijtFdJyo7Tlx5SWwOvTFvrerpphK+O4PW
EFjDZSp3AqX9wbeL+9efK4n/uGEUAHtf0RHh4+WTnSkYPNJIfpBvEDWZ++vCAf6Y9R6x96O8qGKv
kVUMYyonQY3R/b8MejqFg37PWEL0jIjlsn6PCyHvdoCJZIuJfij2BxwHVG0wlSGoZ5KebScmxX8R
xxVtzNI4E29rs1P4I8+D8dMU9pAdr/NI9mOyQa402abn4F/nMtl3vjM3OWQbdBIITPvDM5A1l0Su
Y67eAMnXcI0zBe3GAGrFMdO1HaK6H8ug38McsWa6Xcun/mf4WCQhwezbzEJoZptEKE4wowaNHPXq
FkxSEvMhdXKfnH9qOAw55TBqMMmw3m/R8m8ChcDsEu5QdDIpEK3UAIiToaQG05v9UR+VfYSssh6n
wKpgXtVUE+7MjUlLFueYCBbH9RwzTUDNl2Bw+4FXRqSy7dYE/NFN5r9tmVH3nPiXJJLI2iKYzW0i
pzgDzd96OrCCXCkPbUOKnd2lQ7aKVI5e9prpVs+IxL8Db+Ygk9hMjbpnRrNxX4ArdEZ7iaaVIr4/
ol5tEv55yV+KGYdmGeP4KELHQgUSz8NbpEHrVIY8W7vnV8R+PjnAmdzScF7ejIpB/5nzgxWZ0Iii
0zefrOJZbDSsRpdF/O1bKWxVA0dQ0lbcI1tjgmRUT4pGIWdD08YCRurTC1JdtgxVaNfdxjfVuHUZ
NtgTuyys589ZoPY/kovL2ANoQz2DH8MAgMiXzKG10AnWEbD5xZRLHwSacgzjXjziJCA9evDqbF94
Vfxf9vPnlyaCTYBhAzlMiYb2yoODTlqMyaTdzpZ7pbuZpJIo8WQxM2l10fvhEzU3/mLAYvKIQq5Z
k7EkN7morYssPjkIVA4UWZ2Fb/j7CduXCmImFYNZIlwPWh3Q6NVH65GpCXc6ZFpNhptU1Z5lxhu2
QX9V9KotnAfS/maPOhXTuIEM+NGCNEWr/433CEZAEgbDmEArLXxEO4x1t2bscvr+3uIk9Oj1/Tac
4pnIR0VeD/YGc6MpL0TQ/hbKRaJZ77O7oO24yGaTk+xHkrqTphxq7EaljF6C8mN17Flc/fb9n0w5
adGhmP9N+NI6UKRISMyO0MrT/Ex6HTZulfsmveLlTVr/lRvwnYA9WHayUqO/rtLXMymQKlEwu/S0
OJEPT190228aX4nidXKXYGttPumOagvNiuHVke3myIkgPr3pr2Fp+Spu8ZWmWDUEVqrVTCATerWb
U9DdlLq6H7rlmUHdsdW1aK0KJT+Uz+1U5B8FOBAESphvKKxQIU5yFkKe6yjWmiBuuoAts94ga4JX
KleVMKStoOxo/rJz/xVrLCaiyYWSJWctLs61sOjT0qnG7+jbZu6cBo9u2MgzbB9c+8OlHdXv9X7h
wvLGux6g7WCWtH11e5hX2WNUAB1YrzgTCQP6ovt3ERlV/PItPWAMxJiqllhOaA/bSM9IYa+/oZbh
g9VQU+saOwVZJZoo77uWrjSUqm7ip0KEAsbBAE6pJy+eZej0jqVv9BumDhJ/fRJPQw77MyXjGKPA
OOCPBrf3Tw0mP2ZM8CVdW3Rey7IdbhY3Zjz7wzFcy8c3t7RabUnKQa24S6NeoGaD4go/dCe8KvoN
gfVeWAuYfWTcMLiGk5KMipbyAwiDoYGinDQDccG0OD52hl9JktsMQ/o/NMJalXfiJVCKf7f54Zy0
YJETbVUUwWU+G06MWQ2Le1qvDieHCK8wiWQrgAceQo240yISU+dnqRmbfH49U0mhVFDvrezU657K
eZF2wAfscj52EU+a7VTNh4LdosT1a98hWHrlUfzMwgvZc/dPyGQLlrJkDPxL+av7IUwvVS/w3VL+
IRnV85ANnm4OnAXCFTyW6FCx1VRHcc//5QGyqGfHZR+Kiog49uEAN7pfkQ25aMRpD8cedrz85OUV
yT5FXO/sF74+JWdvDaU5YIrji0DbQ3P27m9F/I8X39Mpv9yNNyfuBtqCasUUnN+pc6/WbWFla/uO
+KCWsO7UVeVjkQmiXYklk5o687TM6kDp5m3/X43Uz+BOlHBLZIMItsTSp/8JiFJbhDV5gEWsj8hY
AFSUFOKVRF8c+U9LrTGl99/n2a3I+9nm2jcybEZZw7GjzOIcGxUucluIs5IixaWOt7VAW7yDPi6o
EhqHDhgt9htfF+InSsFj4bFAVh3LmrBgml1Uoxfv3X9SM2PdEGNY+5vca7ro3qyzxwb21x6w3D07
oyieJDPgJO3T3LeHtUsyL4Ac84+N7nuUCEwvzqOHZADavfInuC1y2qN/PIsEofWMvZsFHFFK0nn9
5thPOtBebJjVxUQSVLLVcJ2fanOPb0vxbYTskCLoqZl4fADZ3nmHANf4eB9vRbgWCZYyvkDOxS2G
5dAK0YGnTdtEAQpASFg6HfxIr8cK+JsnB5p++mTIvGUKhkLEVuI3zM9EpurtnE6j0PfJhIy8vO1Q
b8r8IBnPfKAx8jsaV1PMu0lb6WI12IhlCiHPWD+WUWaLdjnKfDZfU96rhJpy4Xavp5Ii31WR207l
S43BaRz/3czDhIQbW9vTZ4Dz8NsZjvpuJbOTKfgEc+Beez8N297Fo69Ay2Quniu7raXQ/jQzI3Zb
X4xMDkWODJMxBmlUiUReqepJIN63laVKlcJ8Dh44KesyUW8rQGhmx1ZepcNZGt1aYzfvTYdgMAUz
LrrnbcRXP4xiRBTmlbeBAS3sNcsoGCZaURVvtQg147+8TlFEbwf56n0gPczfRrzyNKiCMI5HexZG
ECBHfHTYtN+SrEtqCv1u7dplIXZZMTa4Z7D8BkNF9CVxs2TKNEsF1Y45+GFBCP87He3cAn/cRI4i
KRfae9nEjt5WYpOL4lDr0FQQ5/66oKR/MVgEcePq9mhj4DIGU4oA7cJWt9Zxid061YxE8UsslaC+
iZq4BtjMarW6+54uoVL9Y7DDvF07bTEoF4TmZDNVKNeNMqHcmUUqtFubWlnXn0b+8s6ilUBvfGjv
mr06KDo2/PGCaQgHZqoVvCqRUcK1MPb6IfYeftLhyhRTs9KknTUKiMlQWkR2sj2/bAkYlwGt84JH
xEmtpCS/2hXxjuZVZe+e+xTbK4p29EW4yZdgDhdAYV9S8BmJFElykiyjulnCC+5lmet3moMDYq9+
HtQ1WfM2akvb8cepQDUrsgomHfzHHejeFBvM3SOICzsmrEcjFrsH3Z3+VRNNufZzySymNbqtezLt
Y4wMabQPa6759as1MAxWW9pRn3PZovaA1mc84rVI//zDFazZ555QhhOunWQARK3iMyZfDO/8UyWG
UklhSi3TOidMKvIceyUlGfkRJhKQaOHGwIe7DH1ecMxN17sIdGlZZm+S27nJEkjvfWkFEpZRUN9g
Y2wnjrQQ1s2YbCi5x9QMdMoOX0xRXJqlNMa4rae1vLrFsshHEl43csZYSPBT8lu8+AepKO/6gG0r
mDEPajuYsUz/T3y4qKtruGoTpasaFjTwj/weG3ayoQJaRqRy/gWb3foJO9XDyBvqnejWHeF8ZvVf
58g9BBBubhA19BxzpUaGdfbjPqcOXOhzsOGylQ2GmgK/RtPZCek4UsnPIShnMHYR0kgFHWw3ZPEm
qcMXgxoKDS2QH6fLEg5nykwC8npQVkuoUHlqJJ2nq3fo7b/SocfngO3VmxIMlhhwbyd18LdA2PlZ
/0OpwoCq9jLA1JrCK/4BRzvCgr2rynrHt1l/0AbnpglyWwFUNa15hyaQiksGOvgwPjqPotl/mEjT
FDiHxGhUXSTAHfE9M936PU1Kcno+yRJVdAQUMXieejk3+h8srJvYEyBImrpQqecVmE1XJ2t5l2oX
K4If92yl7to3p6sF5V3SG5OuyQkHNGIYUsjUOcHbphUallYp4Jwcy0NHm02iU21c9f9fuqnfuqZR
+gUTT92KCQsfVpJIa5eoP95q/TER75dcqXd2PezSTyEx57CHMMXJGw+bpL3ypu+Pq2oiC1045wrj
vzHO2jVQGgffVmroGFU5HtQMnLi9GdTkvhV9ZXxw3uXM0EzWZ9sOK8BTfcd36vUpih0utZc1vCPN
bFbxIFrOwKhI2skui2Ds2OZPYlJ6KDmvoS7aumuucnv6vcmy6v3RwwjwRXlfj1QdNNFLV92er/vY
NcENj93NCVRRwcCwC/k+qKs6CivQXMNJS4zj8azMqcdlIYq/tGRpeJoIdubh78mSHwA3uo/EvrBD
jwCOikcm7SbeRRqEeOq1k8CRlTa9+2QT/iYrzYvHBFPn8ZOLvXZikFM7uK9iOVKeCdfosUFdQ9nn
JftGdW1wnpiE3LXjzNpypdU2p4mB1Ea1WvveWkrSnUYqYmNyLmZhxJ7syPAIE5qEWOgmyia3VUTz
oc2CBkjOpUMf4Y+C9uXoWdeafNdl1nSnu7TMojNnTwVA9A8hF7PXFS6Zyfe8aipZQ/xX6cKXhCYc
gH1GVs8HBba/IVOVLZoI+bX750kTMmgpq30u+LIWmxRfaNzzv/fd3wmfQqK1Ph5673C/WYW9DRcv
wpyYUnc5GcYanVXLlmGqLhkWa6PQFcJ6mVoFaOmTYtL3+Y8LC5TRJrm+LCNu6hXeHFQ4/UMXjZfn
QvQtBC1DMpkVQLkimXV0FW3gOm/v4Kwb0S2GfZpOfP64clbQfwn3EiD22yYpSuKSFVd8JcrgkNVM
njUlxzzdls1fkCxX5cJ5JdQjZyV5u6l8MDndadC7pKdZoUJrb6hG9JbnYQfg77do1DsDmfNmKG2D
NhVNXD7cfq8pC3Y37q2Z9yB9BBksZa/uZ3yG2mIe3di7bz2IGXY8aK2mYZ/ABn107Lu07HJe28IR
iAuxOanbcCA3piJl7N8tvKuSoFXtDltuNSTxzcvsT8KVznSueYcjBIwfmmwfHqac+ulfY5VIN2aI
mB+X4V8LkhM192dJeJLy3NACi01CGhwBlITkss/vx59/0Ryk6DhA456jaeAg2FaKzl9rkOc+7pSW
Eteby0x51pi0eVknRmwxUs57hWnrBDq3nzFcygNGUQQgOrcbjFviFcZmg8sHZJ9NosDPtF8+0WoQ
RMgIrufCgoXEFOkz0AI83kKXiNskeVDIL0bLXx7Ht8PkP4HkQtAZRAqSU2a1+CXxpcyAuL3B+/sL
A1Lzpl2sQPncfdSIG5IZieZgFA6jHmqu8urq372m1t4WjlRFtMwRiKLUqXjGhHL9RM4bufyNoc/I
/8fvHzulza9PE+FkpAAs27Of2bkNpy3Rb5xPZxdnyOvZiMZfYLrEXs9m/n9Btr4yliViQ9QIKtFg
UqivaiJ3NQFi/3OqwXDXCDJT6HOaqWTc6Jfms9WN/L7nve5Lfq2VLugDDiC/6eMIhLf1juEgC/u1
cpMqif2Gsy8n9YD6KjXXtIXhwYraZF/Ar2D9weFalH7pC/ppYE0XvwXT7pDzfQMzWMdKAg4m9+jL
wz21VEmANqAocobsbMfFg2OxWFTOqx6miJnykBiQrfzyJn5oGb8tO7KLGYUmTI4Q4/SuBsQz9gU0
LQxdLa8e1YE4sVbOEUWTce8TGkKaYK7vIKvNtd6bLaFrFptl3J6MFOJHAc1Gw8dvocpq+w0vNlOK
sP1kuO4WwiS+IWXnZYMh6IUHfy86ZN7WLRiP25co1WbyWTU+Usf9TJabY4vDq3wP5Xd34UF/r/X+
ahnDQDjlHK9p0YhzQ+ic3Exvot1iU4r3U1ZPLRubBUyi7hTuvzfTr1vgujyMKa9KXVw5EdloGmh3
vJcgMgpvlPNjfChz5yi78M0ZKNcaVcPvvzJvdDYICzyxMoMfdpArnQz4xLO7ZNljdV/RTWiGwI4Q
q0Rp04JaV67B2wJid66pZah+DPR14qr4S2qKTZf/IY9Ink6FfHOo+/viQijs7aUO7BD42GAHbVnf
ICR4xSg2/1cUC3O/cQAYEv3+plwRK4xIWG+tjH4drJb67kR176Ba480HILRds0d4SEj4rX8UjFlU
j/k47UPuVmW6oU+4gEu6xN23eNsy+bMfrh28B73QGbeeoZird5HvV55uspRmUTBXgZBdx9Xi4EiG
+CTDtJNU6yuIvnINVqbcPUSokXcxjKrKI0n6oUWzzgA2qv4oDugNGfHWsdhsdlo9kPK8eVsUF04E
gQk8otty7xv1DCEDB6pkVRTkdM0ZPRs9Ylm++0zC8SjhENM8L4ODH8GL499crDSuduYrZSDb/hVy
JHiXVt8T4v2thHbGE9OV//BahLPBeyDKAj1rEfayr2r/wbvxs6aTgVU36DgxJ6NjNyepLICXJVh9
lQFHEMh64z/nTUfMZOh4O3BS3CKan5xYuFDYb93X4XSk7TNMQGBUjMzTDS5EdlFZ09UzETKrBjGb
JztChqHh4p+NapJef8E/rTDTNFhphhn7ZsLPwvHgPSTEeyGoJ/LfhgRmljl+aCbsm8SlD+yqBRbO
P8YHI0aDk/ctSLL74n97A72AADvC0xUCzZbA/Jul9107baLAMHjF2nZz/HQRff4Eh401bUHGebWo
Cwso4gj+d28qggrvMZLVxRCfLOKKbC4Pn3JSJMAJz3MusHB7TfRdj4QyBdb/gx5KFzehGi66M9U0
EVTep5Sr97nxgc6AGerFwX/Xw/J454TFlNeoql/UhgNqug/KMSc7x1DDP8Mo5JqdUc63kGIB4/W3
7RY/LbcMvSc+pG10CzDVgz2GzggGJ6vqi+qlcL2A5PSIder8EAK+R5kdKgPMhA07sJsJnXHlaruU
L38wI08141CyzdVC+C117cAFN3O7f9AkqP2yGR3231nvg6AAzv09mq7Use1aXVTEwURfaQBB494X
U06U9igdo+4AcQ93YjCihLO5A8Ml8Nkq5+eLnLeEq/jOrhPH0ME6MuOGcyWAAFsd2AOsacztzH3k
bTDgSXiXmhCOGBXx3Z0aiaCDp16yBDUyfODmAK/MjW/9wgBF+J3FipsoY0n3Td97ImC2dRpzkmYj
rq8HtxBNj++8gqWn8TzokhSb91Yl64RKKbRKv3d7dItYSGnsbvrUQMcl/toDHrs5iQOT5clqSorn
mbbFa/6L7uWPnFGgZZGbiq6HE8YItMncRAviV+dKp51rFefNEbVbew1J+FvXfItnRGYpxWs/r6Q7
ScRADCeurf2gsAs/YNXfe7WHT2RYwHa3ku6gTZibl+G5PZUmo1780fcUWY3ebo+KvoaNWBr7tShq
R0JTOE/DRnPMtelzRm8Tsmg+/5SmAUf01JPQ+T7TzOtQrvo7uS7Seu2UjsWhl5tE428HPe+tfPCT
sBDX+NAuJAxFlj2v5DUqbPFJKtfFZl854MXdtBoGgY75frINq93vPAKbOmxWNKpUi+Jmhz3cj4K+
0d6cbz7CaMYH8i57MCgNNBHvl1bfSFlfOpnfKGpIHIa7fZC/E4VqMO0bBhS6lm747ydmZV9SAoHe
geCiITv0xQtVm8C4pEYiUXo80eHbtOAmbhw2amflqDwaG5e7+O33Rer4+Y/QshUSWTx2f5Nb6xDY
82RFMYLVZRY5WVQvjt/q+jW2A9s3fliSfO6TyNA8hjN8JSMeKbTTbIs4L6MzWw6UGgcQ10Q+rTnI
Hq7XzxxjnkZGjRwHQyc4ujsri2YA4AB9XQKW7G0tv9yR23pSn7du4vvjYp6MXLgj8GOwqEM6/lBV
Q89dt9C09kSCKfj4ajC53EURoAWZ5mcFMMlFLw43+R8pVDa5ukMdqmZ/onR3VVZbx/2mMqTDsCVc
NhJThYPfHR66sfDfgMAsrAe5B9wh2ipmedHV1rwmaAQ7H1dOEWGj7Avyx5wiy3jxv1SVGtJPS7VE
5qvQlu6gUAbqni5Q/FETnDS9eUELeb2Sclw9EzFNlOWNpXNA003mo5U2EbqOdHpyrzqKS500TJMd
ltvQ+tTjc5FEgWh2WMMn+dWkINZWpVGdo1BAdIYbmHm/yRpd6DoAJp2/+IBrDUpxjYLCqe6SQmkT
ibg5WtMoO2zV3VfZRAJ8TrocsdbUalIGFXm0hU9Ngqgn2ZATH7kmiBj1dcy6bcIRuKvgqANFWKAH
GrfWkWRQ5sTQ6Xan3gHDJ2ddS63VRoyTKxcs0nlnCY37xGktkZeMclPM7ddMjtBZauYEBLlWZpTY
v+7vDojStMa2OgqjbEcTpAORsgs+pHXg1mYlgiXkRqS0KHWpaV/e5aksMJ7KQkOt4s57H65GO+iL
fNsor/UjAOPkhWSfxRbmGJ2/ube9kaMMTI4mWyz/MdVT7N21QnE5NF035XtT0c/5kqgs+97wk2DR
b2mPibUKPpiLeciWeCUTK8LYirxveCpuf0qcnVckjjBPuSpwsMF4fCGoZniq6jc4HOZgIcRCtj3n
FlkeuQIflu31GOnjmwq30GqZ5K+w115awhUae9tjallf8KPb8IdEs5qv4/5lfIVjbFnlQgs2n7nd
eIoXSA7XCbKj8hZtUiE/MkSOCvOuDZUylCiiUOjP0mJ8X9RsnM8AL765BILKBhPRQSYLN7tm4Nf8
ufSL6f3sWVOVXhKoFvdzvWCdQV1Q7rJgM+vM/+RsjSHvLFKoQ02y7y5VZIivqJqhYtx7xryQmvYc
CgUfh3SxHApd7uqpEOkxRwi5DrhYQq4v6Jx+WhxW1xUvg78ejK+xQBp0X+HraAM/FfAdhb7VteTy
q/TBTlMgHgnc2ipQPOqr8KAo69cQC6I+KdJD+/JvlvNRrIBBCfZxxHpVc2dL5ttDe5q56LUIPvPv
Qgj59q5A9lC98HpP9NNj8Tx/Hx7i3b6NcguMG54djx6TlsLZGKYZU2sQMQWzqmW2pSG+8fNWkg63
zivvA1NnJs8bRnIlpcPRnR21w2qbVDi+c1trGrevKGzboY0TTNtgVXhkzNauyezG86LRipCx4Yyu
h9Rmm97Pgc2UfwJ6YF/8JGELDzrJxAM4i2XNEQq18wFxeLx37JOC1Tc8kxDtZcA/uf8s2VA5l1zb
p6p3MPPKVd2RfZnYXg2IhnCDQc80ruRgE9y+p1oYkK8P4pjichxlSTunz5xxobKyiPq5DQAfdaXU
zYKaFfQops3yloOC3eigZdztBEn9ClsQ7kGZmqCtK5MIMY7yfeldANG3JDwNkMo+K7SNwUePcACD
0qGgPKqs2fRyiuv78kvWXF95tucFwPi74Mcr0oeUO/rPkpho22rehJPJcBBFFFPFk2uPSDWFGCKW
BntrdH7eVq/cLrWI3j/l8F+vQtBGgxIz7Ige2a4+aXjDW5KN+ocJWP0J7aaLAs1qm2vyqP4Pxgi5
GQJvkTlLHcPgwZwnpzgp9lJKCB0TOn5A7komxfgx0wiMibz9Z9PONcoxWRS7tThK9k6ekH5A/LZ1
9o9mxXOHVJeBy2d8/yg+0fo5EZ5XjzQIUT0FxMTtrFsJsaYkU2BT5BiB8BWkyVJuGCmpV/xhddjG
YhaKN1vdeUPemPNdUnag3h1TGR3mKVBveRBHQII2ldRqRyRQ7boHREEx3PzFvVmMSUg9a0em4oIK
ymOCKxX8mWo7O/tWuHh5BTh1PGemSwZDialMwHO0U31N8vlFmWDVPEIorW/CyjwaTZm0ur+z6Lti
UE7l1HYubsEuUUj6Uo5lmXNerp6KuowUdkdXdK2y3U8rFW/XXisUX47hbeTCQJ9eG77hQ3L/d92X
HgULVqXW5YxvGjcqKSiDBovpCF9y3+Gv0KVEQPR4HcoScGiFltCuWFUnbw3mh90/biDA1sWvFUEx
B6en4lF/SYt2qokIJXfnQeapK0hSfLXtSb2rAEZZmrPXvQCeygDvnHG5rTy6cAh5E4zAfYzwbV4D
NnLTrnSISIL3ePjMNYPmkrbgU4Fs0ZR0MGBEfkeMpbvA2rEynILxl+gZQdfyrnA8/DoSx28+6ouC
/z/idolYajHM/0AuORjPQsbCHzUpdPq4FUHebo2N8nG+pp6/tzp1YmFad5xihwM/11xyiFahCiJ2
sj+OakBW/YTcLOE5EeYisKqlahjX+/xkPMOxUXBPL+gWwm2kZhuFqcpvjCLMk2giNvpR36bhckas
5shGJ2y0OpB/4Ptp/O642fJizxe6tEUVT3J79WPUCwPXT/1kLRoa4Z6Ls7lnlo5Fx/AMq2b2cFY1
GGoRtuQIlPv22KfDDarUFn9JIIT2Bz4vPD3S3oktPr+tsoABwlSz8//wX+9TSIFfHZ5UC++jKnSB
UCp+H59sSmBZOoSfqew8Bmvr0RGekiDUXySuIRPavlcT+3UcIIAFgKPbaKwDhN26l5AKo0bWpBJX
prZjzeN13V8invRUASXBIdtId2VaCPD0fDtAeS3XHLi1cBgDw/pa2TVzXwexxSRHEvo+KPh+sbdl
r+yY6ujwnBkHE7fjrEEsdyicwMSHrLYGGfAGTGifLjvHtspU4PuUfPDPfACk9mNW990jT+M2Pppi
q+7zrv8mIX7DZebj5HY2LXvLC5RqQROMBCsgV8koUTcC1mlAYQHMcc+FKm98P6ZwaxlweBrkLZp3
fVEchCzo+HNI+S1GumdjnAlZwuL7Jol9MXC6F7LQ2BI2Wj1PpM9yRL0Apyzhors7GvL3VdeImy5A
m4FlvMoHXhSLP6NednXzpT4B5HDKxunkv92tzoC8OVH114KaI27Etmp+qzLVZ+KB/C7Nz94Y8xA1
XarprTXGddz5rultQys6UPrmaAWWxf6BQMGK9Y6tUw1fGQ6PcvJ4zMrueic9wr/ZAJVtsoAjT7mW
gjUA48qgaR4tswx9BMW8+uoMBioijgceUyQcLH9fbWngkuQ37yxmlK7H7LvanVrGrRen3oDnFzRs
jb2XEuA/bnHnGf19ybs5wyFyL5PMLbhf1p6KgFyRObybTBB5ZtGldOUOaqk5Wx5+B/Z7DsLef4gY
3N1K+lFJoQfgYTY9jcqIf9f5MCAd2KcprQaY0ooRYpFcPAwcXzdIfRZLoZUqRXxq9GlE9K+ugtSt
UUJ81ovMpuADWrHPgMqdi5baWD0bzLBZRz4tEgM7l2EKh7vySaZEGsdxYP/9B7ojqFC7FoJ6N2MS
nzu7Ip6FbKxGPYOahpekJQLyWlHlCcOpRdeX0KYGNMr4Wq42FEJaKJxqV+bdmWtpL1/DWAzGITRx
Sphc5UZdVOicjCnJbkW7O3S/Za3kMGgfyMUOEQDNFLlt7n2lJykk2soqmaM9Qhx9di1h6q83A8xw
artEne2EYSocnMkuVxMBIhplXLKKPqlEvBdwxZRiCXoakObKUkBsP8TSvfuOeD0+qgwpyrMYmIT2
cKkiSmOG5wHTBf/Jf5hlX7Kq+AsNyxlP6NhwTwasBOB2ze2imPa3ILLQ+XmpQ/Bq6HbHP28g5kD5
ZSz4Svl6yjpu+NIc7CEvVpvoahqBMQ8qS3sF2ne1BMu1sTXZnTarFtfDLniFntRXrfYeIgu4ZQAo
6N00kvIHxln+dgwvf8wJdu+trmSJX/cAwfqGzYWHVvk0NhYrmo48MsVcz+7bFKbMD4qX/EjVb3yP
JO4QnwWgS0Bm2uJO82t9o5B9mjtHADzvZFrBYdv81xTNiVuxYFrJKmM64wup6CRs6at1vycCFLs+
ZC8kP24I3lKvaavyRyZV6DFzn6TsVASyebsNrjhcgH0/uhbeOHcZfd1PNmIJwuxFLbaGGL0U83EK
9TzAKXg9sHf/IhLKCCdsun0ZELbbmd38QcXRakS6grP1Z/vd06BXa0tYv4oSIXPdn8UqZBq0DNqM
LGO5nBKmxMoYQzb1dxk9IJ5uVEMQXiYEsH8Dp2QJGgJLfLcvFkvzQ5z2D/zni8UxX8B9JNmh/3pk
JSJDd1654V6Vj2JEHkrHEnTIYipxvzdUWwSnyMaEPoWO0SriZMo1XVhZiZgCX53t6Ybl4DjwQISm
BfqgQPvHXAuv4HXyn93tcr3ZxqkpcMjcEQVnUnDiwsI5wXLw8C7B7JIqbINBvcR/S2M0qmwBY0pz
EvNgyc5ePjbsrtJiLkoQZP4Q+GfXpEiJkiVN74TyeABlOWblxs9gNkbiIP3mK6fcCeRIu388CZnP
8eQDc1W8MWnhg8OOL7L6SUOeH6b+ZzZk9E49BWAEWOGHjVQul/UeAWsVBw8Spu3T16UqsthU8r+0
kdYoy8fE1kiAKhsFG4WkJpTbveWadkDU36zLb+MEZ7um1cBBvrj4iEZqGxGcJ4I6n+mt/EHW4gWi
YYL2la0vxBy6FsDGFSQ0m0EuCNmK13hpiPurhzEcxmmLxj02Vls2p5aSoxwNgZBMX/TtIKlAZWBY
lCOElEk3nSRNY+7OFW+oqivgBqU+msxntDKLu+EPUs2WsMoipT5Z5P8VHith27kg5dkIFxF6pGGL
tlGPX3IqLQ5eFk45n0CmGOJqlXl8BSLfp6ulHzdI1BN8Igb6m1koZnUK+Ws5mCVAbbD1KDy6bk0d
DSnhHAIEwjscs519keJIcmJZ9mOjMZUbYRmRviCj2uRaQoELJ7lMnFBzqP4CX81JpzVkfh8a2gS7
mWS7v9pVmyneydFBxjWrgifAKUnrkxe+XtpAt01H28wFJlBR7rurvUoHdVDwbfMNx7Rz039cbv15
7KOzW1hts/OMeId1E11o4gHZy+ecYP8disjPMPFsB/sat7BvSf/kuQMQXaz4gE9daIbh3+82b5Wq
9uzbXIjuQOsC/bXBIHwGGalE7viFF7xInH5bOF8V8kgoUC72ZJmclCVvEsGK352BjyXS6QZAy1pa
Ssagd3fBlHhQSU79T2RBOUKMwJ4sWcAbtlArrGIoDAXS1D2NNfCweIWJxXjLpKXhfLI0kwRRhtiP
Q+oXCwDTyYClbM/FVkUj2LLRsgQ8DZNsw5l5jhfOAsHYgLV1uN0i27c1cFM6F5KK+IGdVqLGFtpp
ohtFpMdzsvu/1Lq+33I5QttKusSUTq3/t80xh8o4d5fcKR2xLi5ARv/vrcpqWdWcO/25LiwuLq60
bSXYQSCY9BEG6D5Pc/k+pLBaOrspAIzDpcnajsILXClVfSY3SZkcGsC4XAS7kwlE6mzxdTNvY2bY
mZd1PYJ3zOD3esYmAAIFJqbBu+cwjGu22Yef0Yyap7S7wZHffxtbO6UCu2E9xMYjEnogmf9qx7gb
GyIowUJCTPCZpfs8ntxz7N7hFQ/6Y3DI3uhvbzf+1IOXjo8QhOEk32wfo6xgsQnfBNqXx04HVyVq
gnYmyXxue+y6gL9Jdyt9BUyPg+DxJ+wcZabDlQ5apY6U8S37r/BPPFsdbpkzvhXJbzBJqC6ySQNP
EH+K1Een14QXocy+FD+jcISTrw/kePeGjoa/lDv09d85kH6kEckt3dy8onRqiDmCv895/yust8kB
VgLY4cpPI/QADcP0ajS6KYY+qkBfInoT8yBRRdNbG19GhMAERNRUHQahhBjT4Aj7L1nKVp4KnUms
nuWFiQ0nVt8tYDpHXLfRAGlHLz7N9E0JCoUajoqpXD+jKfg8Eelq4lh7pnkc8h++cZx48w7X4+l2
ASHWuemfRB09TSBq53gRNF8Fz9nNcKgVBAP+rJlTHI0rbWVXkGJdy5U1KlMoYY0M+hmbkdCv9n4Y
VuBDFkIghFnVHYIImhLd6UJjUAo1wje4pt5k3l9FKXEzvnnz1HdhKPEWGBEE8i9utRDOMcoIzE0b
XW6cXUnEOOedX80MyMdSvEDoiBHhL/AHECyp1G0PPP9Cv1AwPdrSPB6lzCODAebIgO42WfhedFcI
faN0Tr6b+Xwf/Wapy3In7k/oyTBLxkwljjEaVs8ZziC5iowH7IU6XvFUlOCGmFHe/kO0lty5zBh2
Bd9lDhBC3zLQZwG4clZTXXM59kSRc0S21gn6MFra/ijH5DX8Qj+c5PW6tCoUNN0J4kFJ+1Ks0IES
TTLRqdTuVOXh+e+mCRqPWFhbMuDsv7xz755kyGEFLFpxx4v85hXkGhzTeFr6BtQ8A+8yVIEWs2k2
yCbTqlOE/GAx4+lgb125CPW9I99QzoSG5D30MnoKtSvzFolYuemOUQYoQqx92DGUMg8NLEe4TVHA
sK0syuqR3rCn8W5q29D16CvLFoCPLRC9/A8vH523TiP9Y3M20+dxozfr/dR4rB87UyV+tnOsJGz0
JcCebmqxMX9KViqiXc5UOU59Va39sj/Cdp8W5iWhhXGNiQTqVAvVbhNdQXmn77vxv8n2yv8Dfg0D
/sQ0TJnGQyg7dz3lFAwe+2WWYgqyegOHAWN2qySwymQnz1gNQa75GNakgCWoMRR8XBw+gZeNjf+Q
XiZYZPAN2spgKH4zE17ICEWBW95MBKuWafuDXevs8PA4VD8y5NJJuyIukjX44d/8qt7k/1L03NRV
98r8YpCrv2XN8J4oeneuhANpT5lxk4s77ZBzsWo1c1f+ZsYKHrflaej5iUD3ahDUvohRu8WhWqve
8OBEi4dhHQaJvKDRn7TjjKLTm4kcyybVRSmsnRh7kbuXveEx37Qg+790gQeUCW9H5MFzcwKXI9Bp
hrhOqEMv/t0pWJkIP8Kt0s5d73D3OeeHracgX66GnGoiFzyKwqcwgaQw/CfB/cxOt/Oi9zBhk04R
Pg+KkFBe4yhscNS6TznIN/bYpCN5aWGHNBbi5ggD0ZkbT6J3S6KpqKbRyY4PiJeesZ+1i+5hF3g5
1vXhgO3iEQUS1GCfRSeqpj3lvg5H5+H4kQHj/vrRwcMsn+lKG1jKuqLsdSZWm5VFb7VtcnId97GX
FNJ2+gJcI9kQg/NlGaMSHBpaSlo9ZspU1keJMfDDY11Ea0s/leELvFtyptNtZhCf4rAAHivLK4S/
k21Rsu/ejGVFb385sGkba+nx0z8QOjel5FnUm2Hq4Uu6YVVK1LWa4z1lo+dOVtBSM/FKJ2k/QTyQ
H0lz8mzMmyZxjGyJvylKlgwpEdQHGUeYp0yyuBa6TtpBFA92/sG7A9oSCETSlx36dS6HVhLfIC3Z
IlfveJ68hO8idhxHq8K+pPr98MJNTqz7/7FdazOtYOSPPdIEWkHhrXQIDX3t7+mm3WI99KirAn57
Qc2/91k4YANXbt6JhRo5VFxwhlfwx326/OIPZvChFzuNHWZo/Vwqyk7q2WGU9DamPLfitvfZsYM0
L3pGfU3yTWDwiyS/ltTPgMFfG/5gj6ptMvf2T/lzgQ9l+/Ha/QSyZtIYMpLxRcTkk4GxzuIcPawP
ear7aB3s/PmJjQPdF2Tqq1axdhfDLvj/bCev5Tja0IeMpAMsdyxw6c7Sw4+x6zGSi3dmT2SaK4DV
FR4kI8cyMmLwggVdWGKKmutZ051BRJP/k3hhctvYLz6YtkyPrWSEtiLWa0X6vJ+GOBp1zdw9guea
3qt3grRWVL3cT7JEGOpdzlx2NMslK6N7T5i+7lfXauc2/FcCtviSB4enIV3PSulK3958rDd4Xunu
62rBOLxbqQD0uJnWNXYH1t/v6ofHII5B52KZBhN/oWuaVXoH8QsVf72EvlYxnevAtWTBPnrXWvK2
QkYSVGF/gKKcmzkuWp5lo9Lr2N451Hb8X/ZP0qykaxfGJiTVrBZ0I28P6nnodhSFX1x/N8fQOnQ4
oYpWUB8uJnqi7cFdrULEbPrgAWfpkmh5Kje0xj3mTaYWPC6+IH87jlb3P6PStg6Azn8PPKgwFvEy
LlM9VRqxiK/cWAw035t1MtHcW4wwpLysVUtK0Bc584k/7MhM4gTdot+NKsWEBn2SLfoXjqsWwr3E
TRdQNfLLi6C5gCzQZ3+Chm/I6GzCF0Ou8jeqHbmRnM6MoZtCHusTLfjexXirHi+UBaB7E4YlsOqx
IgtvS4hppJsoSfz1aeqArBAiciMyuZfLInbFDbpz1wHMhN8MxVd6cbF/2XXDMbi8GCk5uu62/+DV
UaPzwuC5SFV00Lloz8wMhe8lXoHvqbT3y0qOG+cPBemifARn9+XmpHd8KSC5JaW3FKf/RSAmsSoh
COb0HGcZ3BtIB27ABz5zQN95YF2jZW/UxN+vKawNlkOihWHEw9n2EuUu1zJuEp8GGiNoxyZj/DDu
hjBiR90y07guYjCXBeJQLEQoOpnnXbXjNjvi5WPiiXlLDjmZo5lFgob7F7nvV+l5vkW8ax4pbKQg
veo+S3EnTM2svm80ps8K3AYNjm+l6Vi57seOQZLUACNkgon7yeapmyXc2QI1bqNC/fdsgboBoVzk
egFmeex7elM73SdM5OC2Lon7zlZATUIBxeM4KAflwgUT6lqIOB//Yre5+7ge+MIkvJ+rVfcDSn3L
XttreO0zUnotzJyBZ1mlSr5w3IvzIk2y/S1dIFtZD9Q9BGXV1BC/ZrohRUGcCA90JSpI9JYNpOYT
Pv+RrB/FSiwSgEnB4TTTVoYq+VNEx3WLgkr7GMZSq8Fl0iqflAEwKEyIf5vt33/gpMcdZtIJficO
gE1YlxPkLXuTtxAXlDYQhRH+A3Nir09AAJvHXLM4x/cwRam26VMNIXsWbEJfEXTeZ69EKU/z9WjY
baCM7uCVvzADsBa3gvjy5dFOmYsnhSPXUvboL8Ij6Ddzf19Ym+X7W9GPmSCeMt6UnDBcm4WSsBTq
P8gao/gj+j9HwzacaHdIYvXN5HJbH81u60HQu0vO6KPyDrqycIUOolfOE0BEY+W/qNT6ZWjxofPF
cnYcH80EwmF26L8mdQqXIV02Z5EPEiks4XJfOzYPDElTNEtckQ5w/OiN353HvlzSZ6pNQoOFI44W
/fw5qZ9PUunWFfkPLXMso1io44G6Drx9wRi/Cq9UrlHJBL3NIbmVHrO2NglT7xdPThrBne16WAuD
IL3My+Zs3Hduul9NVWLtFge66Gob81U1liRedyhqtJAEQx5Kwq6D3xF1b3gl4eFuf/Vro5eXcKU8
znwNbOVd8WG1CYo7vihdaoRr8oRREoo0MAPSnsjLCfLpYVITsHQbOmKItyzemKlSwKB6OH7IUgjH
vE3tp/b1EjlXjx9xll76s+ep7ghQqnzduHT64fc3VdopXyFcIm9sEzp/HM46MfYN3xa0sG+Vxy0b
gwV6vndf+fYVxxPpLMf7ZHlGcbgEgZO2KCIOUVLzqB6xDbTNffVdjbD3tUFiRlD+pNYEVj2oI7r/
c2pkuOsuS8LOR1LMiTwFPxZzD5nGWCJXG9y/kD1/V8uNFpOwWsIXIYlOVX8OwtmU2QrPXZqRpLAR
OTegROJ2L0T0PENSaBnbINJGpjn6kQ6YthK850A9Nj+tId1rRfaLw6ZQdmXRv3kyJl1hQm7C6tpH
PDLp8oPeOewI11xTollLRJu3RdXPxgrfIEi1GfZfzRM+ap7GCNmLbYommnZ2jyH8fYEF/qC1ShOo
F+QI2QBEoQJbtL5rZF3oRcfAgu96LVHr+WOUBX4OeZ134OPNweP05YbtylMkQ+mTWjWVLjbc0Qoy
9QMru/neP0Vgda3PMeZyIMQjCTOmAHrEjEY920ZZex2y2IrwWvCChn9+Ia3qHZo/9Qw/3mGrhr3Z
IJlxDGKp5FJ+fLat9gHsOVdFtyVgnQ8OxyAzGtgemZEcogrhaLdelm6QvRUrWlf5gAtlHA61ilVH
FIFDknD70ZCoU5llgKRR+sg48Jk0A4t3Q7M/Ur/YGrq1O3YHxOykAuHhrxgJRbyMFTDPeCvNhI+Z
pJ546vVHw8CUANCtjx9UZsY7Bx3Fc9A0oTzmiywNe5y5S2ctjRfJHXP43sTDYJ4LsHZX5hS9HE5T
cDCNFxBruYd3lm/Hl1wALWpfbyyHnX+8oXAPbf9O2dhWZND1k5Ic1O2S6LV5drY36Z3cJ+6pIXOG
xmQuOalwIlFdbCLrf2LjrgGBXze3uNrdTXEQh8ZW8hYTpUrbIVKIwRH/Uv2MkFBcoRrQ9Nf0zZ1t
wSY0yxeaXaZEwnfDJODmFm8/bnoyqgACGjnq2ZA6qOBGQaZw54fD4ISIwlKKUHvoImFAOU3BeXIl
K011JPffClGCUG0xecTbPvFfPIjXTKTK5kZHCS65YFjLh4O2VwJ5zyg5EtBfQFSqumWOHiMMI2ui
MT76jLcWx/0Wg7tCSGhfpX0+D7LZ+VcILGoAg6Fbd9s1Cg+ybGp/Wv5o78bnzyXIYjb3bYxjIliP
G7OhUV5KGJUeUyYSqZdLX4XswAGMWzA6wlN4OMEmggCGSfTLRABvBxpJj3oujR/z0/G2PglSbFWX
3tVHEcXEreArQ9d7IGcBEpjk9TZ9nMLtpx3qb3tObMFTmN4cOojMK1zD96ijTAFT7KTr3iuGZA5L
+S9z8QJoPe7NsEJ+XoyDYzk0Zg4GNhllFrH9pM0bUP3XGixnhbUHy9RpHjcoFZOxpoPuUPtj4lwt
6I9kRNsKfzaVXG8L/2QsJmmdRfaXrpP/VL9ESUs+kTvOp1TryHTHfllZeuX+NtA7I4jwIkl6kNCt
EyUs21M+zK3xqlcstQmXq69j3t/Hld5M7vVU26UmT8zpgEtFBBxPYciR6hkohUibuKJCEjiR6ERU
YwZy8w3efeR6YLf6zUBRRITMTFHy5Am3+JToSo4qtU6U+EqQ4EL8LRsCJyapcsVpmAwl6GkOEDXh
gS07hyJWvnXrQbufGH70321IepF6W2t84XdmgaWpsSV2+aCqLl5CP9EBDKCRrIfGa2cZj+8k4Nkt
MJHf5f0VAnT1LBUybyM6hxHpWxzaep57MQmIVKN0qEbNCfUwArFz2+DCZsdC6KJB18Xy+Ke81uJc
4tshfsy8ozm/LpETQe9HgMycbOLrgivDJ/Qu+ZRuTOmSts1dZZZ70grkVbhN/2J2WPw9XYaWhded
u1dR0oee8mFuQT7mpzjW/gU5jrCGzudG2YOVF+ULvbOoMqVpCFjLDRQWD5KCCUsEMENEDzT5C50I
r8giQOkP7J5tvt33lvSs8GuuaDhiLZOmjTDCYhOn+csu29yifN+aP5UcYNZPdv/pglKbFAZiJ28c
SLF584Z6yFGRm5VlIaQTl5bwUilg222D9RwEbGKPrEusNSTcK1sLzZuxn6PJJEHFpAXavft+SKoT
G4pzlY7Mg1L0uBvsqOW7nABpPUZhgU4XEeMkscG3H8NhF6k4ChR2oSuvCZc75VwPqm4s5vR8PbKQ
J5Mpezl77/HUBjpaW2/ts64g2ijZdiX2G0FFAOW/U8WwWM8xg3fKNazcwUvH6dOPceb58Jb+Q+bs
vbBaCMAbIrffTsISMo+IH/BHTzJ1cPtn9lid9uCKjMDcMfczM5U0StU9R+Lemz/hP/SLYlxh9joj
OMq1lEopdsDgpL5oEAYKl5x/4xk0TocpJupZyAyY2yoe2EnDwPJ4IY0nrYHG/Lky0XR9p9IS6B6v
cZnUCM0pzEmR1klhrMoUmYwOR6cOHLcoJvTiUAwHsoXNFUdICe8Vgdval6dsJqcxuKm95hcaWeqY
pJTPNhckpxLTR3RGBPqEyJAoqGwUwnGHhG7uvME2lp4p88uJz1VTphwCYqbc/mECggXcbRVCy2UV
8tRex4O2e2OXynwXteoYBMPC9NMJy4ehAUgACdGs3hcdqXzzjMIEWkTuE1j2/cc0p39BqgL+Jd8e
IsR0wPSKD+/eWXHtOiE4ld2vXePRZTX55CUTKGayXnti7HJABz/axYgEEVsd4lV4hgNbqrOG8nj3
96nYc3UX18PFCYyl9EndF0pWZ22r/Wmc906RKRuixYJI3UmsovXueTkxtjuJAAeOcGomoisWHJdM
gklxnBn7vRVZRI6O3CpC0aB+7MZ+8k+4RIZHyl10jEpgPuaCBKfHz767nroHC74XG0jQM7pttZRA
HFPzdC9euLW6OuivGoV+y6Zjp0G46qmU+TsDtrlfIeG0xLcVmHnolBina0Muvq3/gL1LSbb9jgkB
QHYm01EFyJvv5cYMqHnEQ/QzS+OjIAj8Qy8ksMkceBaG+7GcYy9SQBkDTmBpTLHXSHXFhK0mWtUk
T0LJcFrxmnLq7v+84lSu4LMt30VAIt95G/dRmLiE5aOXU81vm7CO6bIo9OkPH2RuHz8IWx6ucAlp
9UH858sdUp7TNg/69H/xmIAZiys1UkNeyVJoyalvby8jrB8pzjhiUrPBmrsuWk31RV41VO1JmkMS
Zi1M3jjFx+6EMsD4Yr+edkT6kd0erqlYAfAOfEfmsCAi0GEUWvYeavMKitPJr456YfUH+aoJ3An7
E7ZeovmQ2wY/5dpNtYeMKFSGMHecsnDlbFLxvwedlNHrXmbqiMv1hNDqS1wzvL/PTrGwtgH/l6Q3
Vou17Plsx3zQR/C8LbsWOs42mlN/VOFOgTzgMAI/PQII9n1xrGi1srgFEwrztfySuTk+MKblTcyV
EnD+Y1KHBHNupdBxSBzu6N7kZK8ea38V6HyPFKkBvK8RTmrT2nVuqEZ/1EwwU5apFkNNJAm1Qf8O
yyRWi29mSnWPUzPb46Q/hr4zVRLKGw80QAZKifBwQTq2r6q5ZpXXAnV1n01idWF10WyLUgOoIAeQ
U95Tz73g00tO7asgOJpKeRFAXdw7ldmuj4OJsa8hHJZ4ANJyTYfGJMU35Hjh7IAIw2AVLMt06GFJ
uhXWV8kQtvVAQ3sRDmhcoXBcHukfDzfak6OTHnSmiPwn7IZD2HS4uNbyu6BLlvY+vYgb7WAOwcpE
uDssbw/iJIpGmZFTGX6mSsJqAtHBt/Br8SSahqcicAshi8bfNyapbFD5aOq+zgD+jnMa0hjHdOkv
VBnXHErX1vylPME1cvHhgCzWRWmJMxaGzxPBW31nFf+HwFuSyJs18dq7D5iKYEh2lCTsS5UNx7Nk
JqmReunras8wpBq+fCq542doxcgtg/pf9NfErcN7dK6LjMuH0ZOMxgVVp5s4ZHD3KzmGe1hF0VTV
LRlk4Q6gZIxd3nlqKf8rl1fyjXVE4Tbp0J7/u5AbVFOCW6tApFdlSBuAUcAkTlTNNYkHUYZrGc1r
n9bz1nGtlPCSiE01u8FeFW8gsIwkOM6grOb+UQKvhR0r6H7RQspiddLDUXK+46UA4pVgIywZjqmn
JkbNuPMWF/hYN0/Q0VoPDHeIEysGZJctF8Fc/EMwLjnE9blr1TP7N+OfvRrLT8q0TKoxaB1DrSHO
cUHgH1lkxD3XuXmGnXHguPx3/dbDhJeZ8kQEuRVIfp02igzJM95PnBo+8XRnl6rIeSqmibmtYLZG
cdZlA/FQ3OiVruty8NQKfhNV9xiLf8zqJcuhQu3Oiv851NDZZwRGnfIi+HrBAZPEinxPijFyhwKZ
FjGaCBjopR5r0Mm9YTkxdF0tshai6wKTryV5/UDske2UZEoqjPy9r2so/jig/V4mfD8uWPwwPuXr
7CALKRxk61aXREJoe00MAqDmFstwu5FLGrKM3xBWCyqdE/0xAkXpcgMBjhU1+wNRu1EhzKjzRqtr
qFRIvuh6WTtmC3qf3SwIIVhunKHkZvkFICKG2l/nNhFIWHHH50zlVLu0gSmBQR7kj5ji17RB1a++
3TjAtSdYXKnFt21vxbEC9H2PM7t75oUF9NFUc7BPDkB+wIyWs0RGpjfvvO/TGHpIQ7tCtMbO00Ex
TfbwJsGDMG+FnEtflpVtMAa7ZRnQO8kjhzS10ZBlZzlHU39csk9qjychZ/rSD8b83lZaCe6/lZGf
XeVUKUnjCWqJK+TwiTTG6SPW9kDJF1MI9yuFXK+lDqM40ySjMe3/QeheR86bMEkyHjXDly+NDwul
yjlbp7EDXeJilUXEo0TWM5xizujAzg6QsnKzKVh6tgKgrDE4rxnL25MUbTial1lfUkhwP6uuRmJS
5QqLurwQy3bhtwHDqdzy/aDqn8mq2dcrY+bCdblaaN6B/De34FdXs8Dvb2NyQvo5VsPfNr07NLB1
kBbw4RxkKn9I0mP6jd4cYQEPeUCzc3cf+K+21uHnYaHUzm/jiXJy6wCY7aOh8kgoDs3vw6Wixk1u
PVZNB36+QJXvZVo3wRFX+vMphMe6uKLi6HXQjkZqXcl9mIHzBWjR56JurGZs5XW9mEJR3io04DXq
dGWKC4fBCF5uhH9sXJX+1FtPD1tK2Vqb+o3r2VNcUOZqZNn9ny6NARk7wFouTbWeHlFTjT9BgEcY
bJAg5pf3O1fodW7XaQ1bYP+DrmFR19b3bKpN1ZoJoqMZgHTJdyg36lCp3X9Yb6kTGZopfTcFZ46s
8wglenh+bU8qCVvfzOk2pWasWjTLEZGzuMm+xnlTayU52hFtByHph7gc9Z3K5ydK8HTBYV/giKXf
Kj7DSUI6CNEokn3XcF6qhDiJJjHnouFie92TkEvZ8RoIYLaMoXR7l/YhfUmm9xf73ApUbvR3adLM
0JmlvQFCjGOgP8s2i90kZczjCH6W6lNDdeSGj9Sx8fm1+t8paVqArFomBWXBT/7cE0NaamGYKK5F
JLH9YzzDPt23PVzDSUNGKyvE5iazJRum3UMCoHYcJ1GQ3e3Kh7ttnwRnxqkjKAtxj9RxA0HaT2aE
UToh2Gtd2bIqMRUhMZR/W6GhhuborVL2C/ZLpHIO/QtDUnYY4Bg0UVrhI5wdTwcX7HrYigHaxlGS
ikkFRKOUMqqnMfhP5oJag7tGEWJ7iVVsD8xKJOdssbcGm3DY4mO7UTZrOfCptONQo+5SxfyBP7YM
eieN+SkZ3vxxu40ct9FMLC3fFQ+MAvIjjCybIH/WiP9GWZM+cXWfB4JnYYXU2K3JPHBI2K+34BQ7
p4GgSEEeMhPFuHXsDEzKQNrRzfhxBkGP0nvJZ8usI2OdfVMM58krxpmfv3uc3nvEjPjat5foz978
kxzt8huH2VS0bgvA/Y7jge/DN+2iY8RblgxJSlI1gNNMV7flXh39RP0itER6ioXni75GkA2e9r/F
SKkwFp2DnPGnYuDAz5fQ5xWmfkqZ4IxDFZMYOCW6fJ7FQBo7LUnb49u3YQCDLtYdEW13Z9jeNeDp
XllbTnXwv/KOa5JbyH6oOEtZXllgPrQWsSjUIk6XEJIpQkL1FY0GKlrZkuUsVPYOK5gVA7DoRLvh
TuAzOv1e2kWm7r7eLd3H4FYxG3IKQBl36LEHLsvPSqxl07ax2YvBX8KPNbW9B+RRtaNKr4l6fIoW
pM+cnUovfAbOPOaJTFjNhXEgR8cTYE3CkMg8LdfIruZH3QQZ3YHEVXivHO1RYAvDZyGp0FOaqDIf
3cHxFuuI/9wSjlCYDGvr2OAMdlwSGwbb7udqRjuH3Wq4ehQIvWg7FWXaelFmU1TdoSCbarU+vZ3v
zEhrJhGZTCQJTIc+IH9tb+hPAFkszzA/Bppg73qZxMJvgkiv1EOR+3nhot1A+rOGrk04d6DcjMTy
8FpzOQvXlV5GNF6C98vxNdmMd13B0KL3g9skhQ3W7vYp8E+Nox1+BPVvWEXFzFlUK4MKaCVrxQwH
cIu6rGIft2IQFQ7ciEiRh7SPUsPjydBJY/WvBolriFC+T+3uX/zKu0OJuJX0VYwYv9xI/AuvMU9w
7qFghZ3DiF4He8yic2f23t9o7ACRoQiaCrDPSA0SmH4e2q+AZhgK0TYeI8/hU77OJdl/7HS7oIbn
2TLFETM3318Lz0+YrdQJF8UXoYr5N0+ob2RD6cUTUW/Ii927Z8OQTeS7Ubs543xw1JP+Ol1hTyto
M7SQnLHiOx0WCXl+fYnJCUboh/eUNXEIDcVAWSvQk0501NEdISMnW+yJyzZjomoIyYLHDKp6CAWd
58oG1d0bX3tOiKa8i+g10zRi2YCv5LAjITVkNcdwiqyIEi3KVCCCQr2eDwslRSTDO/RKCSq/gaTY
iqtt5Jfwz+lpdBul/cKQSrZ9XqY5/hLMvnCToIfuY4cjiwA61Pd9VjlwTsaff2rCam+Anl7AZY4Q
O1e0rSJxiaUP6Jpoe+GNF+vz7+2qsuMNj3hn2GPjgrWzEUYLCvukyzZnodhFVF37etWxGLiJj8Yp
MY/KXbtDHADyiLUeEN+JAbU7UeXw+riFD4ibKWbMKEvKnjUskVkQgeBuPHwb/kNmylkDox6MQC1a
bneikm+h/liZ5zuD6sOCz+cNdq46q2a6w8KWIHNq8NshjcH709WCRl0nfSqTa49U3TdGRDeHZQxo
0NCyAy6pTKz+E+ZGGms/5dP8SgBOqc08g7Xyyxt5kVKSPGrxpc89DFEo/jkvdn3npGffKytCv4rn
JVohXwPjL2jI2iIz5j8I/80yMP8rtBabNjfM+++XZC7kcFQ4ACPaxCc/1gc7vEQTInyDuQPCuBuA
neLheQ8bwrcQ82apVM/OeAidk45f3Tax/mD8hocstZwn0gdLo+bw8MPEmW43ntQskEgcCg/b2eJS
zc2X5XPeaL+rY5XzrDvodMbtwU/aiC3VUhWhg3/q+7fKzBR3YnEd12Q7WLwJZpQcd4ZHIgA0qsx9
kobXzIqTdv3n/oZoXWjIamFhqFc+AlKFdQrMp4z5F+wogTUW5DRJ06Lid0nFSUwbcUpHS6fBmaQH
KZ3w6JrJDo8scS8sGLcN4S3Gh5xMUsPOpBNb2f0uD5Cqd7w8yEgDPuctgWaXEQtzkUExG61wJZuu
5AMCyrEeDCoF2WC/0XvKBsF6ARw2suppLhuhh+cZF46gahgjqONowTXE1U79wCZRolgRmcdWgoXs
1vsaLUXbUWmsMMtkpWoKxc3Ogb3Z7SDJqy430mWwUNSakF33gcNPwV9u70wJRwCeNNgodVLllQMo
2407YIMOeHKTCxuafdnFbd1QMwPbagobEm3NudeyFiidHoGToztuh1p4+6g00CPx7R0jpZvWcOWg
H0mParqOi9l8IUhbPMtMPAx+QqZLg9kcJxAiI8VWc/ZLeZQii2ggJTb/NPz6a4Ixca9HquI56axR
igcdbSY56HhP+WJeQZ/qGpDQbBDVO4JP8HF33ZwhlOJ+BawOwSio6oxUSRKxJDC+RFbd+RvQq0xE
4aB+VOv+07dYHEKsSKfAa+GlEX6LCRg08bFsX9hdzc+czdWdSa0iyMI/wZW6bYs7/SzgDQNBJV6L
8hw9EbvN/6DCCso2H4EGZZYobLvdgrHFBrxN1Tn+phz4w4lG/bjyv4zFanC3U91lsh2PVgXnTD9O
fcuQcQH5/GVBXDJbI3Q9fBPF1SjxSckTr1JWugGm+OrGCigK8Qr0vdt+xxo82fX4dmufeLDMeZ64
yiMHzmgzjyfiyQLATouQLaYhbgPt2U4kZjDfq8X8a0kidIPmRH6siZWhyG+bsj/eDFo5TYoHosmb
idMSM8YZvx1jbpDOiphZCxoEKD5ubvjWJedChItjM/nh+nu9yZ2zmEvZh+6xn5VujI6J4C5/n++S
4NCXRYz+pSEVkPiqo003EJJMKwp/XLC2+9UndHnQYHk3qkLi4mb6FLsxznuFq/7eGzQ9UvOG2HCg
fhQsxwKr9+86b671TeqUDBdRwnGtByWY3WC+3CwOhBaU2EY8XK99vx0+HvHpOcXIdoLZJPP62zRL
vDcJkI1uBDWgECy6uAAtr6FzBmaJzacNBn5mrcJsz5270oB1n/K2Kg8qxcBajBUL46mBdk9B9Ir7
Wt3k3tBS1DXBteeLazZPxLvKMblyNL0awlvo9c7cea2SDbSaCOizVrosoIjVMM/J4OiKukBrEx2a
F7VfjbbbHU5rfRbygjZMza9NURjlbdaXziLYUzxckZbjqVjgvNNU6wb+gaZ29/GveU6HL63HQFnw
5xrt8l6hsFaI4FQeWTy5tztgW0Gn5LZlYF/7r1BoJD9Oslba9P+cl2pFs1YFaeKSHDAMDxgnMvxR
lfj/lXA8k+xyjZYsUBZ9Qd37XPT3NCv2wbhh6uEd//UoDqQe+x5t6EAoDOWIKFvjE+YA4vl+1dsk
JgnTwMQyUPgHi4l/9udSCpm7QMPN72II81qd6IDhzfmO8mhVgrWUz7ra7zsNxrI6FNC91p4xsIKL
eBBx+tEJvpe6MtX8u3p5BHEyPIDuTAobFQ0r1tYPRbxWPDHZ2GJs6Vnlf8Zd243kb6UDip+vgZ6i
MplEfSLZ7t3ghJ/eJAN/K5o2KxLI/jotm6K9S8niGLIXhgQHTzwIAsXFWiQaG6ubmdnCW/ONLwXS
Iw/mvQcg/sBUBRO7Zl/WCWvhIhhqiZqb7qQ880HiZzzs0UopmcD5F7b3JOEfTzdooCiX13EIi/bq
W1zEgUgdpOCLsYWqWaFM4fbTx+djTh6LJdJCS69XJ8ZBJzsr3CQA8M3mLJ0jaLVk4jMvaekRMp2X
uzGQ7XFA1gXadESxgiN0CiVSIuMANPHUG2ET4oNUw5ntrwDRDatKtfOzGRSDR6zhaVM4I6z4D66F
IL2oc2MT5bocYrTTnWBDFtcptWcrFSyji0EpWbGX+E+golm7/ep6Q54NIKLyIsEJ52epy23e/RVx
G7TPlzoUlaF4Qi9fc1odFdBx0PEG/d7xYbdmaJvQ4SjLLKbtvX2NItiIjCRzAay+Fal2eEymCMXL
TxeI0vfprSyV1iuTWXQqzwr4h079Tga9JpY5kj5Fkz20UvFhI87cXRMVgfcmd5KF3Zs7DxzVNs79
/VLAvxgald/huHGD5WYt0kdD41w8kqoIDC7x46Zo4+Uq+lNO0ZQu2CufQDm+ju/7Hgkydmguh0cM
O6aKKXOsLaDV3eEz6FIiqt/mz25EnPgjDyGUyccCDmmy2qE7v6x07YgwGAMWQ+KUYOw5oUmPwGF8
UDDy1MzT7KiBDsCK/gx9iY7wfS7guPtpYYXfsImqhllPGnTk+rAL88kSDWS11/hGenYRUiRSxqPv
qWpF/tLV0Id9eO0jHaQhe2PR8WSagBWk6aSYAUYSqQzlrJdkmEAykj7agAxQkismYRBEkvN255Bm
iYwmTc9wUegXSA/zO1XWuVuIvFYGKeWiHK4B31KpkFBX1ocL7Un4S7FajZRUSSrxiFgLjSSPGHhn
2RaRQMDET9gkL2I0H8Cx2HAKWXBpRsjbHfJ0Gip0wiLVtRdjWr3k4tPnX8MsaFS1s7NbfIEKyUw1
2o3aq8YRA1SjgWS4n+2L6BY5Gf0hndvQ9V07BAzutdrZPOMCyM8t29g3PEEA5p0e5GriDaDTaPYo
BT51Bo6EmnCqx/djbnGsbK8NEhXjTRVPOKD1DF/GjCYceZuKoZBl5dWY9h3DHLUTDaSRckUF7r1m
XCiLWD7tuz2xy9iG5uQXLJ6JHCaz3L45QA3Jpyix36aIbUn/zOMOHPfUZuN1SigaiSdQOvAxwrFT
XI9wTZqR/GEUsMrqLwEzYer9Br64RFzo0QZdxae0IOacrRJg4CWIHgJgOgSTVSuvxb4wABdjx77h
hMOm88ah1WU4OaD8fg1Di7TZOgHPV4DEDypyQBkV+sD9JIMJ9GJfD90A0eleFt0CmeA1sMjxnNWs
IUoVTViKCPbxB2wnS2UWfPE1RIK78UiFDO3hzIcs7q1toyQF2nNTWDRQBbrDSpoQDVt6AupE1RwA
xgRodbdxX97Q7Vu6TZRN1S2hepWYqYEXUPKkyA1XeSJXl6oEPd69EpzIXcPQQ57gSrIJYdaKTg2Z
cbUOwsvE6fq8i7EzQ8FelxBxxb1Hg98YNVvCAeo7hqwqEmh3d1lGZkpHKsTHMeDVNm2ot4WmDvUO
IiyqYIC9yBRkZY6o9yzs6ff2U05M8nNU7djeHD48gKlbdkCJCeTzdIJFPo+U7ME0aCGD2ybXyNO3
wkR7iWgkfPDHFRzJJY9rB/qzec01uGJOMGKMnW1FK9mUKNzcbR01nEwdfun2lwrgp+wfULndsLQC
HP9SSolY6ERUjgYqUrh1hTSrpk+ATCWhHisWAioFyWO6Tp+fKuG+8yyXIUYWtGgYqHFnUQhQPSH/
NExZSRPhoFBq/AJkVk83Izg6YhmrgLl7B7oyHl9XwGpgy2OMuu6n32+x98aD9onD3xBNNqfdBaR1
FI20vt8SJSq4YVuxpkoMSdxqXLH41b4pYmz1rdWvqpLAjE3cz/OZJUMGxBoxOVRkJkPNoZTRSvJt
wqwvMGWLn3qUEjDFaCkVQ3MdfJub1ETNJgXWXvL/5djuUfdmr84x3bO+Q72llsAX1ON5E5dZiH8i
OxZv53ReBX4MA6jMBxJVfwUwq8b6+1LyjB1QtTFFJcggAwVmnjfqZ8sTfuQOeimkdqYqUzWAebZS
InRmpqmOIuuvkCtS/BRWhsRAV6AYRH9nG+QxELPEIGcpUA/4F6YvANvXowDMuwjIedMgh+Zd+zj2
Z7SIoqjl3lF8Q0CkmOuvh53qoOyqTx57/SK0D5ZFctFClQHcmOarSlsJZT0/e2eWQba5w6uk4+KN
G9Cvb8jGUu87EMAeX5Vow5p3lMvvkPrFR+bvljyottt2j51S2xolL7sGUTyOdjBSBBHtwLxZ8jXQ
28N94ANMOmSODz3ww0zPUUGdV4ukPtQTHqD0RePPZy/oFKnMP3Zhcscb5l2hmbIvm3pgIUog4pHr
APcav4/gW2aHEbTAYgWQTsfXsWFHKLkTlC2m+4W04xHEyqR0eFVcOL4lrRF4kpAGD9XhtFYSdQVh
WX9Uz06EWzIzW+pQKJEUtBkGJiXBXfwUeznaZAK5HZf3Wry8xzBU3u2UKjk5wiqJvlxPLvNspLak
izzDLrk6ptClpdxiuC+OV7PuM5wb88Ip238mO/qcsA+7QQrTVhsF/INdKK0Ns+fqRAt22N2hjpin
K/inG+57MYadrl0M+LcWnwC78InXKYu8WTqp7/3z1EuwQIdYSC+nOBGoE0YH1uQbBz6kO4DKNnh7
t/UQZ3wLvgpx/BkVtiDYn9ktxPHBG3wARQqZj/iiNMJMQbZzJYOStEd/GFD9bLsN4SRNTVO0LDO0
BptiWqZ0chIVk2mlSsZB964XhzJrSE6lio+nX9j7Rwdj+6xmkIXuOLdDzM6kIkSo/dQDaZc1e8vl
RuW7ouolDnDSaAq+SpZZ8tJyvDLSqtnfzlVSmEQEcekqpGwFxyxW0zoitD25syVdgOOjIyHlAprN
0+b/HH8XtlND4ryRxUz3uf0ua3WVxnJPDJbQbleZFh5EGVB7DVi1H9k2WTtVKz8y4VGwvViCgHhr
z5wBbEuWv3RCN2eR3kX/oIZUUNgCwL5xYCCmBGHYevs8567u6qjq5OPRP2BnVw9rMBxQiN7jYs9H
eCVB/DFdlA7nM3YKb3PJvr0etpHdkRKuwzCHrpIUXFBiItckOp6zJ8TX2Ua87Ro7s8L/F5RrCkAJ
SNxbGL6hxC/aaJsXUHOSy4wcq2jgd5JATr2wmsJ81SVSrwUHnW6Yp/5E1DWN1xF7WvVlUa31x+Dt
65D2WoJVL2/mx6caaEc85yX7VMB2E4ABv+1f4n2Cn6hKPfDuKIC2+EfmD6gtLCjZDC3k9XRQAaut
Ne7ZicMyQ1X5WzXJvZQk33OfyJpXaVPqDj52rXaXFhl0YBFjpXpIZUQHkMX9kEbJO2N0Od0rS/wg
MfzIWicmXIoMKILqYs11DrdPDf/4iTO+fSzqTpn/gThNumN+vXWHr1wxaj2UO72XGsdy1FHyOpwu
LlUfNN74vPlZeWBtGfsP+1D6sNbWwEoWOmK05U/uAnoWhjjQGeYfp1GQyvSUT5a+ezZG88bwnozF
QmHogF4zgA7uoWL8TgaTRhsXkUdeadodbJ58BOgROSKn7hBLeCcn8QGCcP4W/PT4dz6visH8hSX2
zHBck38EKAfUAZPK3kleyDASnZEGPl6hXOXtQVSi8X/Vqip44YhV2/V/AzHYKjbgI3mExrjzqqFe
7Sh99mrDzhOveZhB8A01xsq4mF0rKK4EAQFjT/uvobWSXsaHmmAUoDtwGIehFwosgaCymhmuQqGW
zpC19ra04NYTn+7zFpZ9TBTXZNZ+94WwZM+JhbdTpBfAdituRryorNbsL26Hv0uAGMJBP4FAARvB
PaRbX+NoxybXtjliXKykCOu8s6DOMeID0iIVKvNEpfzfvLzMtS8yT8qBNVYEWTSzO+w7L1wnyJp8
xvUk+K5cgOf1W0Eikj7NJH5pdd4qVL0R5EISdB7k/fWFmoKnNeXXf3DQ/L0vrogXWsMYZ4bX43fg
EzbXjD4vUQMfwxYSVe/CnaEfYkcvb7SdceU22vvQ0yij6PU0SVGmqoa9lPwMjCZBE68PG4y3KFm7
uReIEzFKhE4rKNwcku+KdknNJKs8Jz6jVC47RYIRYk7sOHj19vY0TLb6sjej/kXE+MvVgleHpFb8
cHhOpUfxoyb9BCqhoFfxzR2D5hV0fFb7HiVEMXH1w6Di08xJABC/r7SdI/05TFUoUVRozO6HheBo
bvcmV2r1SMrjEcG6xEW3mn3K2o0pLCnV47Doyk298tRjVEq2sJrWir9A/tsY72n/xva525EgPMrM
QNOkshmc+Y4LNU5mIJmg88PINt7ZasROTAfzvY2Zupj2KX4OmMKEmn0F4g1Wq+Qa30wxwzJdbuCw
YpuU4oF3VaroZkEwM4Qin+pq7BSTsfgpUSxUMfFZ871iOobNJOta+HJ9byv2x8DccmVH3A/2bQNa
V9FufVcHVoVGPKYv7s6x3j6ELpyKxcqIMkDGCqFPqnkl9AK+Ezi4lGhqv1fu9UpqK+gCXaTxovx6
VDf6Yj/AhCNKxnYViNhxFEvAuS4sxXDUrTb95rhB3YMPAoC8S6xtGpk/8XU7bRxsnaHgOcfCyp4v
0NfpPLXdivx7YIVRLPTkSb005oWTe1AAEka1W0p+W50n/kR+FgYCjlGfwUYfEXhbCtqvkHsYmGhn
NiljO+DFpKA2+sjtHK9xDIZyaq6dKe09ni3hyldkh87O7FE/LsAtWBQmdL1rHRbRBFLwWSxnHY3A
sYTmDGh3CIlxQwULlVlmxLA8SNrAzD6Ee3EEByg3Mvitf5EFEXTeKCbDZ7XgeXB8Ooh7GEKTGMtG
0km1fXA6dfTJnMy1/E09zKeuXnlEwsWg0SptJ4Je0vF8gzc/+EdUYVd8qgNV5yZBPYKTPx9Qw+OB
ZZwdgzdutWhN6xGQkTofBg2cgQ8K2NnELO+XVwQ6o+A7b6WCnb1+sckZuIMDsRLc8s9uBfOx/uuk
H6JFu47bjcZfoJtEqPTGLGnbkb7DJEA5vyZ/60lFScgaviylk73Luoc0uWAHD+78/j1LFPOdd5W9
ySe/DoBWWGjvtCtht1cqAM2Yz82jDhFkDAvT8jmEfcNkOcsbtArtuyvKPP2NFNh5rMZyuwsgUWWR
NaekOyDtAPQ580nhPV7xUElSjN9UxOCgiPqP6ex2Y0WjzYU5k3Yi3YvTtSdLaN+c9wBirwG+x5vj
hYOF6vSB1D/IlMQE5qUNie7SpMTbzGfU5AHLJQSc1D5Oucy+ntbBZJohQtxAEyX7J5rqGH0eDrkl
/uk7KB7L7YGrMNs9DTOi5DZfgk6YfDHcSvOTzjBX/AOLcG9MdLTvj7KkbpI8+CVxFHTott0cNwCZ
f97Zv9xtVFVbSId12ZlYqBlwffKwOPJmhB82GEUpMeL4Q1MB5ISjuYOWOJphJcZJTRjpbLNBKgvF
3Bucxavs5IrnQTO5WjO7TW8yUxYl22YpHUscYDNmIxMr4RrRYjDpBBdypmDYFuxAt49V+BWhMots
XJpl3VqeQY4gnKMvdSmDLjzWm4aSG+7WWQHEcyaTPrkJjo8QQWLtZQXNicv4XraquznioukfCjpN
jSXIlKBnWsapk1exNZaaSshqDJXVSo22Yl6/SKMRNUl2qJJQ7jjX9wZTXlv6N9tIl6b3hrwv3PPu
eWI/BANm2IbkN6T2xP5qQz6zUhyAQNHjzbjMRS0/nAbYx0UJ0BgZ4ongE1LpzuLIn1tFgtWNnuHH
O+AcR7G4ttST0kiwDQV33slxXIKU3vmGiTYhc+ICKsVEITgwJCwpywlh93YnXQQ2fFHsab4z2JUo
6TA6uKnYSHuNumiOYkXRgTbctXP3RgsmO/VrjeDeVdrpV7KxMSiw5QPDvOzmbaQtc1TlFeBl3nXj
D4j4P1RHEgJvD3rDC5STqV0diJ5rqQ2omQAYeoOFnQBuDcgTMd0/16dj/THfubJfqjFw4Stp98VB
4kjfR/I/UxlOuy76jiy8q6NDKnGXQSOFn/W7F4sXtbp0bi3rbcZIw0rAdBSpFim6Zq9vUCo8WGj8
OwZ/TvYHvUs6HJOqT1wr5Ic3eHNciX1m+CmM0lP7Uik8zMnS5V93cvUyrZWRJeJzY0kNOAIE5RU+
7BL6GS+BTYHW27+CbWYir1GBuw8mpyUP5cCLpvF7OesT9IC9E/IrcOZTq6QMyFyqhvqc4UuO7dsM
P5eM8Eek2kWP7CyZk5uS3Eu1KRtrSMsJzh8rwaSzr8wU93RY2pcYRLGdSWOJY9TuymMKXLIgVJZx
Dq3kzY2fxRIGIGKTyknOR7g6xAf4blNZ3BhLBp7ttb0xBLPlhRSQKAkWZLTzXVzBGbZ91cMJm3N1
OYSNzQIy4ptOwM75kpOmNXr5sjohWUTAgXTUSEwc6mNruJZOARDtlJOwNgJp76eqe9CYezE0S8V0
lTWVapc4YdkZ4paRyYEy0PzCVcRSESdpvq4kOSIl7Uv7aC7f6G1LFOYvmH+fRikTvFAuN2BnsBuj
s4Crezz/1lfBOuYGM13QpYzNuOvTzfxehk3Y403Y9Pz1qjS2K0cFpLoMZxC+e092long0NNtpyWp
xNRcatZjzmjCR6Z1SXKJkmsNdyXSW1VCgVC5gLecAPnsqnveAiyYM/MWKP5ehX3L6vHd2d+4znR2
uRMuDD7XeM44oGoS8qJCH4miVghhKICYlo/JzsqLuePMLoStdjCTGsU5DN7nVRp4pVD0UVcGNGH/
MsV8hHRfTcKGJ242hTMM7/WqjPd7ahxGPSTi+9/7Mtqjbj5h9u+a4ih613xREZPv3Fok/8i4BAH5
CBXl5b1vPBVKuYvbyImJ4xRNVdE+F2Vzv8NL7T8P54mf4ZFbtKfTsbDyOD25U05Miley2LhPAuEo
2guxXYELekfmCLdWvx/s30urG93u7lC1h01EZXAdapOCmBRWRyFBcVnjewZwxOlHOcGxbOzxILOk
Om6n+W28hyezQOh+d9/Yi2dyAzoG9zYBUACBjW1JsVATBcEcLKH5Tqe/aZRYU2IIG2pyJ3nhuiAm
4xI9iHPwoWRlVVff+nK1mN3JC5AGrzpaSjwxYtieHz6qCxo8fH8SMCiqltrrKOjvGr6m35JTzc4w
/eBQUwESQfbUVvdYJxokLxiIbBu8SxDcmft7ENxyEbfy9QUXzz0ZglLgxljVG32b/zmEIVZQi+s5
8aGnC0VkInzT4xJorNkcZgObcgecp4QjrnntRzRX4t4FwCR4H08bqRx43/MNzdkID3DKUlqpjb0Y
n4qf1edkvFjbwbZM8Rw1HzzVitIUUX1Oqq8s2V19NeyEweR/GGcJWLUjPusKL839WMtVgBTxGBrb
4FMY4etNnvqmj808afsvWtbJDrqb6UCR5U43HKl3nnWP4pk2yT0l3X7iBBrnzcNuxwlVjnZ+J9z+
7sbE+UdZZr7hnYoKWrU+cpfhWy+2T2vhd8E627CS8GqlC27QxdYUNU/LeqptoJBH7UYHZSpPBWdb
qmfrUONo6MLu1kQ51HUIdBuKCVSSeQm9IwTme2XoQYpX/uLOIaXAX8T3jbG79D8KK13FRry52GwE
jPProwiVcjJ8qQ/3bVDv3LV/Aff0J33Kg9Pa4Hskd9htjNzKhnBXAKHg4JzL2jsgJfDC7Ub2r3ZI
ynjy/7qGe8xz7YwgBibR4mSDbI4AKsX6ClVHNBBkdBckmIZqizIdwzPkQ6MFgCWf9LCNvrGdGGAG
Q8OVA72fSs1kOkY5mzEo9SgSVzMtGz9B7WBktEwQFNjsddsLwuF686kPn141136HzkoWMRMvXLaU
C+LR/XMHzs8iJ6q51inUHTevdQcZWjolBq4DiQclYboy74WIqerSN8r49Ni8Qar3PEp+3+QnRwYv
+fxbEKu+XfIFodVNzurNfOb1wfITe6hvuO1+I/Pbd+1H/VzhM1VJj7nnj2MCv6rCQF9g0UPNYvJn
a/C+UWYPZsUgFfpbOxSukVkGlELqFGUu4ZufAwziycJPuVO4JL9zrCyYWQuX+PKMNftkuDNiQjek
NJYUGhI2CoU+Mmf4XHxVYqrewot9yTQm7+2cFcY3RvRrkHHcxgsz6TvC2xLEcq5V0zznTAKjJH9A
OAWmcUWlh7mMXWlBMda38L/ANo6EkkzTDrvKilGvMPRYwGQcjurWbRb5hUxL+2M1gkunMdGEvReD
F7CcCGn+FfGaOTkDLMNhzlyWMnvwvSJ66azSj9SbJ3NQ1V74M4eugj6WWCy6pexZMJ1VV12Q1IGx
0hpcUrdmcmVdgMMP4pEp+oahDbnyEbDa+VwDi4m1cEk/T9z1dKP6l0tFzXCO5nG1x559sgbawo3K
BlXnUBNq3KmEIDYAUIjGbGWkRBGnsGH0P/nAdnQgvFTKC5cnve2Nj1agB97rIOo/eOVOTjNbu3Wb
75XOnwIqWoWGkf4cQZkaQhPKfbf4YtO4bUoWOQMRWxaFZBvJVgunRQDqc0rS5+8dbzMG3xXl1Qgf
Zgk/FMfcSiAkt615Vx5wovYnUMJbN7uFNFx/6MLsxqi6WxtnYRwUkF4+NuwDkdWgla3ipTQyWji4
2l8NsVwOLRj4VzOe5mw+TZmB8crvcDadtmGtC6nB6j/jzn2jBc2n7kXQc3sX+/n+vuYe5p2uIhvT
CDKX+fCa08+D88NhGQTXDfQtSt4ZMj42Z/FkbXqlpdZZb6JXUkuXzhvelBc02prImtnt29CobnoU
QlRjJ9gip8J+t5RAdFyQZPvDnBLAxDJh8nRFQIL89miPqqKGTWnUV/gjL1KG102uXbHYk6Poa8ne
uReKlGHZc4tLGyLu1MG+tkPElEdGwtuBHQxtCpMmvZWydzllf602NsjCDLYP/sUYbD5RrOBNOl0o
XxFMggq05DPpfO6HIIeTo429515YlJUJQLClyX4ypKYOHRQyEb9IF8DVoaWLzB2Mn7rzwNnQkCRy
Zib0b21KDfH9gjzO6yGW0hZuouxf2OK7zvFelxhCyvlXNXGMtLxmuxbjuOq+G7d6x1L5p0zIItWy
KA1+Az4Pl84u0Vs9D3SqwhCUfne5PKi1i2lsPLpGGqjzXW77V6LuZ6Y+WF+w8NmZJoedh5myKj7i
lOSOTOzFIG1qI15/wCvFAkl2EZvXD//bScPUH22Iq3f3y0DAUPKLmqSfD88izFZI5e+98fUm9xJz
LhotHQ1QwGCB9xLodYdmQNM1cA05dSY4FgEyyW0ZLW5yPlH288Lp7K2BOp+xdDyLpliabM7Uh7V6
VpgCAH4jWF0PDrprvhq94SU28DPIjCq2EBpcCjxpvfiL5LAZzb2uChqz9+wkRUrvnSEA6l32FRfN
mSgQB+xlUqzdnXkuIAgUeWqo7F8HFitdlnnkV/DAmwRCT3B/7SRbkWcV60OCsLV+d5VtbnSRHdWG
MzEmK8DG4LMdgqqJrASMvP1euaI8ZAAtvHmzAB7WjTUgEZidd11IY9ymRw65y+rUxdSyA4nblAoG
UjK+3lZQ8zewktP1oW0o2zT4TCKAW98IsZijoTBQ/mb5PJ8nUDKEivorPqubNOF/UJZXKe8B4HUh
oD6JjL4U2bMcsh5EMRIoRKSHlYeMsk4XPtMakj9SLOb5JD+35Rrhtj5EPRT3z5Fo1PG9S4rqeab0
NoPST6qmhNFoAQOS9bGWzrSCd0y/BdHogzO/1CGWQvcDSEsOqjMlAO0KDLUahUOTnBOEvgScyi/I
v0J/ezEfCChzfxDLIJIVIecenEB7n8qeRvPdkhcRUHg8L/vkFRgHrIhADQVSDbVOgMpd4275uZLf
uDCZ0rYqMnUxyYMEBQTtfzlclC5OQNK99n2F/PwIDegh/0dbKkALoH4sHeK0WoWR8VkxnHM8mDRt
V9KwfMRoPyAOEQHcN5isimwKervxpqEJlB0Rpjc4ecRB3yzx4S9f9jhwDbhNtiCvwib2LYVJlbl0
hJZzCLhdbIE3UIfccQ8Xllw1JeKs8DTrOrDqGCYRKGZNzf8JOZJqakOzis57Fc08/DU+GK0qf0C8
yeXDM2zBLAvx7uzMGYembwmB1dDbP+0YvposXxaMLA/Z1lWJezZrrOqnjsxmEnZA/zBiqW8l1bPE
aCtPaQJhlAyzBCp7vJFwkjLtUoNKbB1SZiMwiUCDix2rvbVzJ3x2rki4e4ubPkRMHHywU9Vj8clM
u9iPN1RoiGWIsEXhV/AW4/vJpOsCE1t/DKdNF98ouwgVUNeBKOykfL49KzGihh8RSelUDhF9uIlY
Y2ees/Bm4C4IzyhylILmNUwX0rlSQDXxyfFLoCNFSEtkELAWjODbMrAINEgLqxycifWWA3LH2HVh
QNcX2J4o/CxkuraGoKc8fkvkLbDbiHxxxWTfU9M7N9PIU9FSkVC/cV+TamTSh9SDloQXbJBeV/Tu
njVK6ZtxenrhVAmlYg13BMxN2J+DJqJH02Jsm3OXrsv8fgfBVwtx7wPSLKsdO7eflSFh8B1lyq+c
szxZRrzgCTIOvduA6Fi8lmXi4IrSSWa2WVS4z7WSCK5uM0W9DIOqAvfRdPIQ4Oy7mM/D/OZuGsvu
c0qhuLHfmoSSee8GrVieqWT0QKAiOiGPUnRlDkA0c5Y0PLUg6o3p4frMp0UDFCCinmDnjGZxk0J9
lZYrfvZKufb+N+FmWlPeE6y0sEjSFMWfKY+hddDa3F69R7CCSh+RvJhAk9M3eWYpiGt/i99ldfdr
fdugc+2MH1mE76T0OKfFGd+5CAlkgQWVJrrE7ItOHI5qLqhQ4/jYXx/RYSNechkHu3Hsk8/QkZiG
jU8n3YR3ctmgeTtIe/4VhAt3w+kIi7FyvF8d2KVwd6ZyO+31m3tykBgnB3jZ+x9OSk5b+ekJG6j3
ElM814ttmwhel8F8xGoONp4k/q7drO24GikC4mBoy1CWySkhJowyY+J9c0rD65g1LAOoy7p+MO0r
HnL5kvyldRDUrEMh1yBLjQ6WGzcEufDH6MOxdXYJTwSBRalcMisNB1zxlL3TYZlBYempLR7CT7+V
C7V6LR9mayOMMq1zR0qEGZEH8lDywfa1+7o2NDkxsXzab/3HaSh2TUIc4hMWXYcXX2M07rhjCmrJ
ycpxWLC7FPv6ncEv3JN1gceo+Zvqwo/1VWScuIfd6j1mPqndRq8cKfa8fdR2+PtuYi68kX7U4HIl
jxC2DwSuaRW3hH3ScME9VmegLvumGxm7hIdKNYqmQBr/avDgRptn81JRyTKVFPC33Gm+sDhAfs6n
14CD+NnYhhcFXgRtH+6kFmlXWc4zdGs+Aw5lgHmJdBEfnJBTpP7FLwz/JIeDQZXZ6VBl0lugORWs
LxiW12Yvzq8sX4CUsPfJo1GlfYCHnjZLVNqrO5UraOIPYkZ2bpVtreAdEIgHbvaZuq3mvVOKhQ+l
YCdzdDgyL4dTwi+DD1659yfXUrstXj7jcDVTvDLHJu2Z9T63ofOFzmTeIqnSVuQ5jfIrABuL3JPM
NDpl/ugYnYrGmwUn4Jj9UcOk8sYIFt0qLy8C8Ynv1z9NStOM8YqBr2EZRuEnwROUEH82YLMPuwbw
Eqwc3VHv11c/dIfwR1GoNhSzqpK2Mc81QQVcJSdzXiT9dMibVslNf8ljYTSg/5mc+7lSTyJmuk1B
jV9j72V64kWYl8lx2BScpJ3bAny/nvLSr1jRfUsOUF+17MsjyWJU82O3gbAeT+teNXy3wmFX4BGk
sQKySVjazJ9ddM91vtlKxrLuuKOoA4SOSdGo7zLE0af/e/7vIFzGO0Q59GxLqfj3sfvwmrleuif/
Uy26o91CHX5e0tnoBMilOK/hqg3WoIH4p1Tb9pUJtxbg+1dKeU675DsLAnuOSDbr/NuutVCQKA7l
/zQ2r7FA5L+bhMygdV/1OZx8CEUGc4GnGVrMXCq2F0HeS9nCyjh3gehxYTqlAfZ77TIUGaSRibr8
nWUMEiRMh5kEtP4b5ClmBIhmZsMk1DT2nfZVnpVvWs1scBYnE1jNiimZrHyw+ffpJyJuIU4YGMcx
6dBpvo1AP6cOuksciL7dN6BmWBvTAEAnomyKNbbc9NxpBLiQYoYCpOnyVumhAhCmkM4osi6SNdUV
qpXjcZVDPZSHGYyHoyH+GsMRRo1wQygt+E3SBPDy9kAQVn/TVOiioAsZEMohwukRDqW7brfnPXeC
xgp8Za1r9ZVGVKOWrdgWsY/gCXK8OZA7aaNRo9HmlAXj2zg3udfdg1GEDNziSNf0h0ytjh7MwxDF
UvRDbXLMjQZO1YdpFJv2toc+/tmBGq32uqTTjItoD0sNeWBkWJlU2M+jaez6OLcQIjLBk3RYoWoy
vX1AhowhQUATyrhF/GHltlEo3UFyj4tGok2Nx3PsNmOLfz8lgZw+imYPI4q9yVBm3CZV88JMI/1f
qf7Hjfd5HoN5eTueOc0QMow22Tf63LHRZKZ2zue1fdrEVjR4QQXFk9idlNI+PT3SkdEKjWfpUC6T
3uZN4esMXdLYwk9vlnCUnRNmi6HW5ZVk45mfF/kp7uM2R6okZFPYnTGSs8y8b9cPdyq68uJOtHxo
seChkVCsy6yrfdXr2X240pEqq0bNxlGGDH37G61xqg9/OBKFNxbylevHau2HeOkJ3yuZ+LIOi1kq
biFuo68Vwc3do0xQes/0sztb/KBNEbhlP0CWbgIE41tFDMunLz+CvYGWGLqQdov1gmMJ153/p51a
DyI4kGXofNBIrogz4UkMFZQteDepb9imwjI3E7toM7sjvBObVc07fMqnJ5fsu9m3TXNULyojrYru
R4Z1byMan53M/n7VnrL0r967DhoczVWsG9viiTX3D7uO6zfiiSDfw3J7tXjXByWV2lUvMJZGIMHT
RWVizX+/ork7dgdVS4QHyfGPO7MXVLkPZLLRBG5fKnb6hpKlSQirtu51tTlGG71u+24sUm/nxYcS
3CNhEYu8GjdpGkCMD8XkHJY2YnfrmKsZr7gX+c05aEPR3Txne1X4ldgqpFMRtYeKR/7jECjqaRcm
RLcH+8fl9yrdx7oS7kpc+fsp59Dh24sSB7520JZtPij1uF/FTQnLZkTaub+kWr6lj+o55cMqWq/d
lZMUhlRYWbBvy0Fb9Y1NdseU2+w3HYc+TJUDmreYfWp9wLOaYbz3lE8x4L49sFODqE6rjBMf3QLE
b4gIiWmV66XYtYTdztQfA806ovseTB1Af+8r/ZxzKZQqWtBSl6V0KfywufwhxTaCZAyhf+qgjlFi
GPWsR8zKMrq7463C2YQEltST8gUogmxtTi7kU0f/F7O43/nrHiIPBF5amhE5xm6HODkG4YVVKCKQ
Bwy7ENwb4vsZvVTD5tYD1eLHlnyWZj+xgxUUXgI4rTio5436K4w0r8dv37YlZ41i9VIfJzLEudjd
TR/ZQnlku7aDfGi2a5nNCm8B8Mo/PvQK+9L6wUTNhq50Sy+OTPkNab/6FwBPX6H3ZBnJvxDW7sF9
lcsvf1adMs0d5TvdX/TbAa77O92zo9hzqRcYWeIzFkliqYEhr84CeuS4UvJeXei5FRU8SS7i3HCa
lwzWaizatBYn7StJ5zbm2nsVANgguXWKXV7ggPJP+sDB1L8uTNORRBTMYoCpMhGGt0dQDGZZwTky
e9cHcKvCsn+kN+jOyMgG68A5XYvR7NSeOjjX4zs+CH+P5iaOCKdscMEyiaNgT7OXmSPbDNXad7i+
29dGibYibGkHlJ/c8l2Db7sPtbX1+OWtwdN3pE1aGZLanloyZ/VYNWs1+cbSS+WLktw3nykiUZsB
fXpBlULqe/82OD0SPiUppJzSrxt0gWUg3i5sBzjghxZnETwmc9KEM3GKIbMVASOjHrCf0w0TolS+
xrjKE/Yecia8g8nLqcUiT8B5M4ol6RMYZacIJPTf9u6LY4lAiI8BeH6KB632NcXvwnxl+BKrDk5d
xnb1ikDU7Wj1QPmH3c8L7FIVqcrYcMYejhbVOmgaZOGYeWejplqCxc9GX5+kSWP002Dmqo/+8e8s
MC+UJqywuXlrgryPxP1Mfo4IW1+/tBUg8QExgBFRHsXbwIEViUYws7RzeeXFNfK0s5IPNF3RlDSz
AH0e663zYSy7aRKcdH8CfhCiyjY3V9SvKrLPq78BnUXDwVJiqdzGVtGxkR6aD/pc9hz8FabVcutX
eCAgKR9LTEhkDGOoYj95M8p0T6NZLEcgFkAEIckYbOOFK7APy0CvDYV/smwA7pdLsQUi6QZsp/Ev
iMDqIYIKajQ4cleufNz7jqdW15pCX9J+34S4Inqm96ibU4TSC8VeWQjwN9/qepxwNqVkLtLIDQC0
ALdosxKis9Fexjrm2gchvMj83F60j3pKMRkWitu3DhY4I1xh5Tl4P/4uDMrvFJAwmBQV7x2wwTDC
CBfqRzhmXNP+FBxPi4vg06gpLB09iY1Gxfn4YG0G6zCvltooZi41BJ9Q3Rde+UylH0WE4w04Emih
7z64Ck+5lQfZMsh9fDLWeSEjU45JnDNIq8LbU4oEDGqHaIrZcNRrhmifutzKZkGcCk77Robzci/j
LxLtdpabzOf90zH6hc8o1YpLPgYMInVGOuFEBntwxtoeZYJlj818bNsLqENyE7In7/8xMxWMPdQV
FBTOvCIX2hTKRDn8osTmM652GbsIOHaEShefAWF1nqevCe54m1Vi8D27U2SUjijPtPi95ufVtFY5
rCxuQLCsyEVX385xuBJimMfbQZTSxaCFVN16otFbkZFslxF3lp2iNOdTdl4yqf6wOheBBVuHhNjE
3jenG+0lKf6zpn6bv51sPauXU2ZJI09be/DrChOVd6n3NHvBHLOCISJ8yRRzDUoogqv+YaIrIP12
J0nBnLXS9poryQ+BeyT5aR6q620mDuaZB4++yg87na/2SBvFAqxcyJyNopAR19rnDZ2SXjg713L2
i2+1Whms2R59wpf6a+plfaID4fzNlcUGSWIwTWiR9u4Ma3gIvr1GByn8SfnhPA1sQ61SR13qSIqz
/msfzZgwKfE9PwpNBro/lDqXm8tRh0aRuMH8BhcS/A6au4IuAZDmFQpjdgdMZDBtGHisiNXQq+HK
7sS9f2YzQZmGMXZ0oAmh1SBWuUZi7i6paSyawQf/nNN4/MOX6vDKUq5oggQ3bHnkTg30Ty2IqrFv
/Btr+e/Ux/VxaeJTYZcs1luCn2cMiD7t7IxDBHd3XWYyu8TxmqjX+p4wC1YQwIyqHGxAGfNU/u3h
VpKPQN2A/iIdi9yly8hBT+kQqdbm84LXGS+WEfHIFoeJAuxj30+5Pe1B4TX56XGzgJp7NB4t8x2/
5snwRyjr2qOufdcyRzCFojb8dYqIF/VVWpgG/VZmn8Xv1sVNiqryIEzvmhb3FBoYzYcmvDGLtfdU
ukvwRkT4Q/eLZAFLKbpGvEvjR6FjfKLXFQaJAnA98wdN7weL6f8w2QPwbZLpAKZaafXoGg0QgvrY
WlsoK6D4EGQU2CRoG0mKY4F4P6umcaNyWDxP9ndt7QGDmVwQ4HOnD0CRIgSkwmGW3lmWImi7ARWu
D6K6dD4DpxsEN7MfGuzKsiMRUq1Ny9AWnbfTBexDArEOUcn4JP9eg0A3bLZ6dkm4avfuFRkgIp5y
4UL5BkfmrokxDBTTkkNKmIKN+mWckpHpg6b8iuGhXKNn5LhVMLgY3bL+7YmTd+d56ZYuAz9aHBLQ
ISfGoP9N+R0fk0WlQ0rixAg9zw0J8EE7BSeSXL67J9I+7OMXPmoyhnJ/EwE0nIIs0XzRZIeJXmzZ
nmRyqgxVFcqMocplebHCd+gLU39MtTkNWzccSgHDU1NopPhAnfkSLOmuzZfZYz1SzcAwcZYj2gSL
ucenQ3/YspDyW7bv2r+r+uii/sv/gb7Nch/N4mo3g/5DQbiQjJM+G9LkyFb7kBTnh5AQDyOQq4ge
gj458/mxm57jLty9++EADRZooOOQakL+9U/UD5ICRMlCldP6bfJjsj5FLRmrds+HjmEYizwNTo5O
OIUtK/1gorooT9Sko1SIIyrggKps5iNskJLQYUMSx7aHveExOT2DxLTEwJN1cEtiR/bES3eSnI4s
2xZ6pJZF7MJFPvt4lVCcAvT/g1r7Q45u1sAljPfrOw2DbWn/R2MJ3RpE+MN063PWMWIbXeodIJuB
P0PVaJaa9xpJOs57f/6wkYRdUEhORut2q8uaULmw2pQU1TXmC8H+W/8TMECZzCRcabqAnRB1wg50
htJGqWJUPoatHo8yuhrFCokMKvY++IsboxKkfLZWL89q4iHxXa5yUvG2XgwO+ZVBEZWXm4R4WLVZ
7SIOBigEQl8DSJADhNellK84lncFiaAwNueZNMGTUcO9KU+wbEYvg+PIDbiuv6eOZ1nU1xFfZ5Nr
lGogWpVdMq6cBq0/NnZZmWjqjRxn8D1K/9kkSPVpLXL7y8NWGbkpQ+xWrtQRTU9RLJRJQa8KdT+a
yIJHkIz2ki59nKu2s1RPUJJI38X7HTlxjdr2eu4HqR/Z5a9lCZgsNELmyUYmH19Xy+ZLmaHprxxO
tpFWFx4wt76+P0HDmH5RcNJrQzBKebrZNCkfOynDHo2C0FYqJVcvX6bUyEpoQbrWpV6y4NYwzTNL
jmHnODCeHeZvjvLMxj/pkRh736vs8xo6ZS+PmSyIbX7acFNv9WRywaGJ7C0E7owFkExg2J8/Ud61
X2hwblgYen8ddrpLJ5Qy6yyJoEplFMvdb/fhjFFH9LufGg5GTSSnQ6gil1fimOV+HToxNbmeqMX/
24q/G1G6eR5qqVRb/MgRGSLerD3MgXC0aVr7veOzYimMsocC2bPEpL/KES0Y77i2aqQjzj8MJZ58
JJyGmsaExGc/ljwJtGVAz/44FqhZH6chD0E2m8+z0gHaubb2vC9DbLZvEaJe7HlDApSSzrYJ/JZc
mVhxu4qZbESUP0x6lCm4OFN+XzdwJUHn6XFlmI/jNR5C7qpUiJA2m3u1LpBRojSd7/y4vPck9sWO
J8HhhKR6MswRboapgs9P+b4BQNJ0JkpPhPwlAS53OlGsJLcxzfBGVx8lkxmNnmPW4B7LgcshLmJz
QCox7dxgvTb/Nfzm6TAFpnAIDsSkTKDGHn/YRBrU2onHEPrHkSF+BC6WVh3S1yR3qZEEaGH8J/My
zMEnLuZ1xB1WHSGlEryr7zpHwMPYcIxEI2avczoJAZP8GzNrgCCwJ7GkYtBSpdKu9QvOYKseVBXw
ry9Dn5gzn7yAs/UX5vWmX58iMHQ6+6o/8T3PVjonnBfAJhS9c4mGVZCDXBBleIP9LhWz3w1FVmWL
MH5ZIiuPX6tniy0nZs+KNuiCUxsQPM+CRhKyWBwheJIU88ZzI16+9dkjHrxoI1LmoRXCnK62Pe8N
ALhri57pnVBF+0LAzgj6WZkNb5gZwc0sP15Vdm0Al5AiuKh3lC4g1/sHgYkKyQb1TEMZvGVcfd0c
fprFbl1Isu8/Gj9hje1lUkm7HRDkkyurcTKWrSwwvEDAJdO/C/5b90k6biLtoE4u7GoYp90FIkNf
Y0yAf172cJ2Xc9+4EEgdFTjH3ZH/ji8aFSEo9F1vN54HYpLydsBlkjqXD1yf5e3F+Xs60VBaoeRy
dRhP4lpJNBETTr2fQ6uHMkXOCzufgsYfhgfMPpmMNrTB5S34gS5cHqBDqmssIU07K2UeHq88qjGC
JTlQK4c9xH8j1be43MzrKjWmeZXV0biJ6CPVTI1XlRTAMV5ysmvxnmcOgpYC14HVu2LicXu5MHf+
+IyeBQIM+rlpo1vAtOIc99bZ3fL3A6agkpBbxxkrehAjz/Avk1e6ZZ1bHHrKLtMxl+FQSu0ArAKZ
77Fv3VJ1tgfpW9C6f0AdlR/5SVxR+TqyqdzG42EY/U7qTu11dbGZeCInKaALgFRHmkJD3V0XgW0j
qoFlMmZ6+YQp+/0glLXTSCuCkvh2BKhumTMqj7JsI6h/ZJiTc33i7FAe0HwsgUh/uC1fjwnWlGOQ
taYJLsCxH/3znhF74QcBXjF6L7lZyYExp4ABpDSg5oIc5NmYbYdWunopksWdQ7afFwHP6e5oeY1g
rR2cEaOGEUfBGCPqvqUHNg/QcjJmFeYhFVg/zj0CDDJqZLPpBrsTSORBMhuoB/n51lb+8Jh1BMvH
5PEZchCd6I48fdyLxusJJBT7ev34R/p+RMHnWWx1TeYUBZZv9THr62BBQwAlnrgoDIuHuBTqLgfZ
UlDhJ2ekezZmwEOEOl/mliMzREdoozMMtG8uHNGIGS/FkYIb+H0JhFjdkwi4HexLFWmmsBPjtMPy
6XwGVTm+vePuaMWT04tO3gU9ERz3RKUkRYIso0ByHVB3dLJj6lkP4wnKnQJytWrCudX5lmqIg3rQ
6m/dfXLI280lUKid6dWUUsQB0BW+p7bGwHGr0WlczGNg8ujqfcg/ArBOMb+k6eOx9UC6jhO6wwNp
M3s+tAC++7RTt6zIYl3NHTTdEsYkrSeBjVgS2/omJ1IvUVTY16O4WBfb7yYF3G4fiFYaeC/rser2
FhDyckT2wvMZmx3IPcphUyIUX4Ur3sdbRa2RN8SvjF96FctiyM8Gbs5FHX71glTUmgxn4kZZYWyW
L/LKQHCzzVlvls+2MTtfx5utBwtGW0fd1OzSgXYF3S8FO6Dz6qPvNPJin/k8aDk5XJ8I9Pl6U3RE
CkMYKi3440vcS5i1BXi7HtrnR2sLlXyQeObzH/Xiqsg01APGAYfcbtRrszFbz6ccxaqA3M4ucCaL
xcyn2G3LpJSNrdmcTTUICUbPnmOjmy009JAwsYVtUypvPly55U+F0ROlfDNT9YZcj1jNTMu5ZoF3
qaQ783d9deG2Y4ZydDkzxXRHQajIOvzUI245KQ4QtLuzJTJ09P8KVvOZDCYOrPmsVBYTvueZ/ymZ
7uwI0DbV2gvj/9Gay/yDiOXiMI13m4/okZ2uA99LUDJ9xNZLkV+AlvXB8JTPyThdYRSljup/EmzT
ej1thB35GJaZi/WONnlM5c+fDgCyJO9Dls2GSfHzHf0ZcYVipDNS/Ww/ijLtvyxkLfQxCaBT5dlG
pebZTxLdFk+8vZTnoGTZHzR+eF8vPYHAQkX6QlRaHZqo1jwYJeo72tqhobG3/CDsFqaYGq/r0e43
sX2UE2iK+f2k1cywKjMayE4YdV5AsOsG2eEEQzRmmYtNtK3P7F//uAholCiVfvrYxSYIb37DzRpk
suy0QF0ViKC1qBwOfx0kGfWMwpimRu5wVJFZdSpn7UZk5KcNqh9ZaElLxROn/ItfJ5H+wGOzdbDC
HQllO4ohPePjUF1JXjK+9XAgvrGzkdxBcKEPuN/nwZHVw9uUeO2HGSeyaOzhoeVBxxFu8b36ofvJ
ZHgg0DnJwDa5VJtobco+eVir7WLZEltidTnkKHz3Ady67N/7C6ThYdaQvHUqdbOMB1I/8z8e7X45
pl66FwT58NaHamuOTojVzMxXNkKKDzdgOrTWO+AL3CpFLUFPCOfpyllyNGOCW3KKjN6xSww9gYM8
LiN+37C2zaNv77oZclQ166Bb/JtXwwPLSZgxHdfCYNFIE9bFoe1+YFk8IzhEbo0QOp3uU4zJU6Ck
n4qtIEDqPSZX0eTW8NuGcRSkKw8PlDVVfEokyEqiYltvwIhFOcDnf+1Bp+gBoHaoNN777nCTtogW
OESG4XbdAez0emwlq6zvARADkc5Iv087Pton0+OEAVqhFvjuAZ7EuBb6jYE2TkJWw3aJXr6eGi23
B0Oqeali0BOtUAGZBaHHAvObQBbYGCHq4n2jKOZsZekfnAyIY33Y+4w0ippAMqcuoNrpCQTqvXRY
2i4vdjNpWs6DkQ8XApH0hHgHGYmX3hqpticyprRuA5uvJm5gYkLkwoWXGzGbqWCvtTlMA9u+YkEL
8YX4m3ehQJFogHOg0UCa8jGlYJBb3ithE6nt/E4UB7Sh30tZwQXJGp3NiuzoLmSIaqatDDmNfhqV
zjx51dg4lqrXIttnVAERpfpbmEjrnc/Xnz1/0xBudo7Owya57ODVi2ZQXkqS1qVuGdS+mlmuDALf
ZEDp8y7I4WB6XJe/VjNNARTXvdy148bgDJ29swXxlBNxlXUuFSpGf2DUPvMfMC3MmEDxrBLv76uL
cl7nBycL+SL1djuBs70WfAsQFaVRAaoMzpxZmq9bLoADr5MB5ZCbSf7WNLzHtdlqx/AM+Am4WBKQ
XpzMYBld0jrUH49/mlh1vpKkHUWL9AWJOjeTtQKi5iKOOmxHwxjvhZSloXxWTP3Yv1MEZsHKN9U1
7EqplMC8v1a8BT4kfHFpt0C+qJPyNqgh0j2y+0BbiVTCxtyoubbsshTRpUJqcFVK3LKqdgWLRkgt
WnYzkye8yssH3RWN7PQ4yXHzC0b4I9KyBWz/xe3eL4iHs+SmHxqeuY2nRdAv7WPrELR7Xi2jc8HL
2TICCulytZ577AHrzoJPqEJFAvCK+8fhghEgWvq02GV+ZEWeyFZ3kXHIdMEHEDbrfBJVWlwm7ruh
KBAdShitOzXy0Js+min6JQZJiLPRsJC00LAIg2P5q42Y90ys49SsAXt0+MG9EXmMVbK0SKW3Unq3
pKa1mFHJtysbRc3PjieGr6vlu5CsZezS/yyx8mbqr8+K52Q8QgQ8UMgzESJwTZxUlgxtaYv+g+ev
KA+GTME8ZYnr7Mct9G8h7g/wmEGGduLp57h9KZzRFcskAXe9rUEIEmGvbVgDZX5es9KJ6jKNOWp+
Z9p5S0n3BcmDspNs4LmRitUr3QkmiS7Aru4ZM/flIq6Hmv3ktqzyVeSUC4HmKr1ylR8nSH9IxqUa
zQIEbdca+UOQYAiIhSaCZR8HT8imgLTyEoHe4XQ75iSRrLhDgWifGNbdhwgszyqUqBLWDBoYtB3H
Bu2K2Y6lebROWl86ADgxupyv5UtcUfvGunLEStfJ93gjYldzkt8WccQtk6c81Ml90qlvp/S9/SKi
FEGUUUzoydOTH8Cph0ViVbmcHOxW5Zh7OxgTR2JFf8/Kuh+S0t+9V2yHTef6Mr8fbzcZtN950fTU
wHzUVWs9uHMfvr8gs+LGKz7qoZaweYjiCPxRQXWYZDs7lW+msEtUKNer4opWO2cP/6CGlpt+nZPg
ScPXhEqYQPPmbV6FK+h7cS8gF7qhIU/kCceAJw478uFuhkzz1SQdpvM9e4mVHpVZry1M8SeRquRw
vbW6YyU9sqRIQ3T26Q6Fa0pU17sGE2jdqAwsJflbFYri0LkIX6TPu6m2tC8H6BR+a6UfR6NOCk/w
Wr7YLTTsVzxt4+pY/cCZ/YXdIgyq4BnA332EwKLW1kfZQA+X9f/vprgacLsA70RTGaOCp7WP/VDr
jLg+5xNdfvhuV2Bgl3qVYKtGQSYP5HU2EjxRFl+jZ2h3xOOH9LiuguHzSPZioL2JywrohVwWtDmE
1wJfBnnUXTYfvjCVYpUHb55oE9JMRUCsY4Nw8ghPMxav3daAS8vGDn+doNLGty0lKq6xyzM2RsWb
C0zZPNnkCfTM/P63k20cZ8yMmOrEKXS0MXyQ836VbFcz004+kY0iJwOeo6HT7l/JlC5QiFw/lrfo
fUQtBXrupJuhA12a9LLRkRQtpec7yAWNHbunR57MREUOfQvXxehpvKMlZBgEAaJgngVjU9yDYD1V
ji1lbhFOkn9FLhWojvmxul5NqVPaTAZw8UOuiOLgfkT7H2oYIKFViCGO+VtUka+dkrLk79r/yFLn
RAVrueqsoDr0tJh/UPLiKljap9Jy3basxkJqT3ZKg7fjHHZM7E3OmBva2awz84VXuBtLLpCiMbJS
nLEKxw4YOjk5QjbqAUEh+rp/VEpWChADeVycZHyi9XAFwRG5ANz2Rmhn92DuYMWAqDjJMMa8HXU7
hwnKhEKZv7024Y4KP46kOS4n2766iefRw7FtL6Fwm6LZ3zLmhuwkJ6t/yh6pRM5QxyDyOgY2ksR+
Uzt4ntpwFX3hfJ8rX3Tjvjqm+mpq4pD7AUqrHBVIXM5GBF29avggBokec6El7kQGzyq02j2dpOhn
CKjXwZwDugKlLWYHx6UkgVvPhp/3GdbaHls78sOfrkxcvuH+6YPm2BMZGt0uy0VCMEhxfSA54zcY
z1EjHKu1aqXrCkwlZPrG6Z5aMkSGSzRoGF8ZyHyDwjRcdelGsA3CfId/ZVFgSaCvpjdeXxfSM17B
Ap7qfQJDx66B2yORROPtQ5Yuqg8+GWtrKxJyGY968S0SwILdNZbFgRalkVRhiczCraIGzptK9LKe
+3IDhKnJ10ZloDmphDUIY0zvgLygzV345yV5PTQW8aQTKXROtZyy3Tk1SuZwiEyfD88ETjh4VcWs
7uO5BAyOtxCexRwMIkOO/oV7aICExRuRUI7KH5MC21KMZ8upTVl4xUEVL84FPW42Rhf2fxFEbYsU
vB0I8tPKHebM+Cp2DQzVQcBOQN1G1s1djX9lH3Q10Q05xbFl3pS7vZ9DWnts5fCCx0e5QgyP2DC+
yY8VIQgFvd4bAaBc3+5htolmlv4IGHYFlEiTXH0irhi9EoVwsyjatnw5yxU/aKXIvJ1qfQ/E6/Ie
xByGD4rAo04A4L/MfOk0NoxLVeB8IC79Pk4urY5Dp8yjDXSdHR2Vr75AdojKN4mKQUVbq0l8XfyB
wlPEtIpKmQCaujOy6j5hrakemaBUHUnFfxG1HPp1vjPL9l7RKQy6iuBNYuglijJtMopbDhHuFDI9
u8n82urhmwVuvlVTSV1ARSI8+Puo8bqgs2Z9ELPj5LbjXCA79zCwfDBp+KNZYlfiyiO8YYgtt7Ed
MQGbYxn0S2F2CCkMSIhfgtegiRLAXo6FRo0LRNIImq2y+4fniw54vlvgMIX96fEeuY49ffQ01Zn2
Fx16vvIrf5ZjvRyZxGR/Q/47k7+MAsyHnbWQNiyH6wJXpgqN9EhX9nsYdNFDOOZaba6Qd/AiHBXz
HVxR3paTfYwtprRZvxRlVr7ePMO2f1HBN92vgf2o8OZhJl4+B2472n6xlmFMNJOdDH9WHkabqNN3
yQz2rgFgLJ0RiuIvUj+awi/oZrGv14yD6bTpY7vkGP4NzE3EEGzesRC46CjndY4cYI2ebfekCfuo
+qrN7dDGn19xZ6rftlwdxgm6/Jw4whlbL2vtE2oJrIosf4Eq76qrZ64kgiirl6VE6v+cm6xgeAdJ
bufbfXU/m5icdfmqnESswR1Q9x18H5CVtmGPtvIsUVW0m64LNt4EJM6bmFBNcTFVT+nEIDK9Ky7x
DfS3S2KKK6wl3ZolWXfrpVLJiHI7rjEcmBNQkaXO2AnHxBz8U2/yh7opji2HDNQYSYEaF2FtmF5q
q0AaehwykjclN5rTcrIKskp6Fo6KrteWXvvtb0enQzjZhQ+o0lzWFA8z2SNvFZ5oLESFh39ON/r1
EkQKDdwKRI5/d9Z/dByuXf5jmYVwrVzJGrcwl4P06AQDtJxWcsGcvnq8jAp2bQpAC6Uy3Ag+DU4b
P4dQx6ugOrZy+z5PDmyM3aaCz9vdMpQMTNn5bSmBaOXrHmM9i8pmT82IYANgXP4VsgsAUSxW77kq
HWD/wOZuCAZNouob0IPGJaD6fd0SUwqpd0xe8AeWvum/GpDTT2m2ysDA47heY4ITPkvZr6qbVCUX
nwOpOTJYnjg0Gd4zpPnEOpGihHY+7aWyDOyCqYU6USnI8BEoYlH3PgdMKqvjSMxBe9mCPwZ9Xw1F
cdoAlGwBUqXrUipgrqYbEC2P7ARIXUhikEhID+2QmiZ6u+PWC77+R1848HRy0hica4dJQ1mM5RjO
om7K8HAybenHtrpJka4wC3Wkn9QFLaVOg2EKiHq89FCWKXYoMGAao9YlA7YI2wp1wfC8QrfqLMid
K4WcmKN6Qyh04c48nLn6RNOfvi01XkdERyHYGN6A3VmeQl4xi3EaQdp2DeD1iCeSLfiYNW7LX+KX
3xChDVRMgHyAsJc6/Whd8B+PN65z/4upmBtCGfT/UsZtlgrsUd2c8lFrVSVRHouD0KT3ON8xGkXr
nLSI8hTng4A4bN9kiSsOjogNWCSHQfinTA+YOQ7pTWzFIrfQ/+lFzdHiCwURICafxP3qJGJYfW7y
d6+Ug9JGfSVllzBbKKjD4/Ni4KZM4TPhmdaCHBgeP+Q2fFM5yyHHUwBLoHVfoI3aBQwBvhqH5Dhz
llq3rJH64C0m8Fz72gIBfpjjjyX8D4bbYKb5sM5bqmH330h+pv0lktSmULb6yzrhGeoq2rAcQVPa
3//aINGWbP0YK5p6kp+jgoaQCmfeCZIUoBYn4E2NaYK2UiueUn4YkDR2GEjuPDQn+1XFMyxHIo7+
vWJRCswZ0TFRKME2jqFsdsjs2YTaKa8j48WsaUNc/Zz9oIawopz2u7F/4548BdW+jQuicmBz/hu9
qqwRwSyCGI7lLTUAR1qSpOrkhDNXvHUqhTWHlmhut6Gc0MDkmWQH5YC1jjMLexxZmtmPlokRI+m6
EmOnoLS9IIbCucdOoMakp17yYBkRf8IjTUadeP6X5Q47e+kqFDh5frGx+7Ojm4hz/Mv1HeUeW2tu
WYUgjVHbIMbObSqJcRhcdpbPefvk3pTTWN8fa5qh1D7IyEtQvfW+Y9Beg95Zl5GLfnlWCpCo6sHz
DUGq3TGA2133GNLqA90y1dK64Det4Qmd0CJO3gcl1BFbzLFx8/BoQDMBLDBd51v7AnH3oduQF//s
+4ofQ4AVmU65y0FzxNANg/Q6HQwTbFEXzI/oKaVcTaSQZzpmHvd91w+PB+WoAd18Lpg1UwvjNZtH
DTtrv6CezR3blBmaYBlyer6tzXT9fjyA8pwkUUz+0jJ4VDGmYKJwDTRTqAc59Bhc2LZqcqkQdaKU
Bd3BlUkzAIrnDcj6Bw4XBI8f3iVVaxTz/Z8OpIsEabFkhgERQmYb+NldOzcfx9MwQEp/5Da980f4
LCsEZLTfZ4zYFt87dphbPOOx1dPTSAMmPucVSZjbsKEG6WiWIkxFxHrfs85cgsl939MXg2fF1HA+
l2SfU6FyDzmU1XrTJylF5oSbjFE6xCTgrmC/PeEesJFco45P90CDwMjD6XIUpqvmVla9lxA+8/YI
W+W/tU6G6saP6klJiYe2TpiZejNwbqKpF+8drlmLySMnTOFHPnRhWSpYCicFZiDUfm76kU2f7qDS
S9wf5MCOFm01xYp47SUVXQoVrOgp6VtC0gS8wHII6IkJOmXHnZJMSnmZn+3cBe0VHHtUaAtjqo5S
AYra2k2C4B93E5yPh/PDBcrDocFqrtSiatwAQ/RKMVMHbpTBKEsd59CCwUxES/ds5jR4J1SfN5qh
aTkhRv6MBvcBKX0ja49UWJI3CX29TZ8OQVBO4o0OmuRg0ynn7EdDLqeta1DaYYPDEdeMPSw1RUDX
RXifSsVZe3kdi/f6cm+fcjpdXvBORrdgtdAzWnWArQ+STk+UvZUJ5dYvAUa3VBq9D/MdG2djDVNQ
2Z6H7nVrFUsonTpE88nYLuelZE1dp88G1nkO0WogHT9VPsucw17xUbT1z6TXLL1RSDKaR8+szhdV
006Q9Nix0iTAbZbPlU5qh4NsVGucsSkUYGTckoRCTYR3rwFmfDzy5v/Xt/2hNRWBM2FQVj1Y86BT
82Q/mbr7++05/zRkenIxlEnsNilrdWEPPPNFcoF2OsxHyxB+K8uzRv2ihZErMa7Sj0/bER5T1rFV
HB93YREVxjCJMqbli7Zs/2GmTOukCcWTAkxR7SF89eQdgHibhboyOR5B6VMFzuA8lb2C+CdnMZ6Y
GAErudjcytvw6JVSIXjAP1cZrYuqdnTjKW/24nLvJ3E9Dwjpc0aaTKmgMwbOpvFKknGq3xNvAkrt
xywtIgl2SXFaoDdxSu+G8tOFjKTrBWN7B4FK8NBmxxngwpq1WyZDcsUHHmeq4FJh9dp+4PAIc9nd
xeS102MMKlwGSQKFfTXNqtyOLtewUwnFcXeTNFADaSQsMxxhXbGAAxw5g72lG6xFYwmFFSr5G2u4
VLI0pf+NDPWjtEdNNipu/OfCrCTFgRHjFted0EVOGE46SIgyoKTbSe64vhnk9nFb3xIYXd/pN0xH
hBxumpwV5gzBRYIxUWX62bnWtn0vGthGWzMQORJ8GeXIgYytYIY+T72OUCfpmIUGzg/5pwDJ1Vts
NtppC0ZkxmWgj56vqhPKKm++XzANzHCcyMnHWFeLCS6PkwxsHSNn6Kr6Fi2Ej7BUgbScKSHh3yDD
rEyPwfKVRffskKZVS2VBcONB/rgdKgkheW55qpnsPxiN7sM6M9ZXgi3WrfOYLlZ/TOT7QN5xusrG
F8dicR7J7aDg0qDQwnHBu8Lfs8KKCg7HI0mKP2VGsLqFVSNWXJDF94gRmsaHhHT/cI3j4grDM0ZT
Y19ANtAgeSiUk/bv4hFa/8VGe59vni43LZZ+6dHbkQMgmLlr8Xt6GEEFCgQ0y3XT7LNnOUDNIi/q
mddIRk7Td3hVhR9keHwC8fu7SDU2x2Uy7ahPuOlw/DThtV9HtmbMW5NQ+fiGS1CDTRXf6MkwtqTl
ybv+VC4MpFc4+pn38wO8ibVFu9PEZa/s31Oc5eNjWRzpzpphQHgGxrE4Jpy20kO17pnt+THg5lKa
ImmaPzpM2mp60s6u3m2p1iSDIKJwUHDLrsoMw7CgtqxtgooxfML4OzUr72a5x8BDiRvNsAbiGjmG
a8JuWugh9idQNu8vTcIurBrBNTmmsaKd6FJgcCHCF+VT8NQx1FmSolWtpCIgID+mDCww9Xwc8NFp
rPH+WBVtoIAGJ+4mn71NgU/1uGTS4RfRv9CR7y8NE7b5H0zHpAgzJ33dFk/ImjijbbU3hosj4STs
6G9G2W1m7Rgj+kH/xBApj+5GFZ/LgVmu6fM6MOwDQvZ7zzwXVwdp2fHoW5d0SSNpG9KO6jz7KP7a
XNsgvEEu3IZDdGINbSySb0PmL3m8SqVQSYDNbyvfkq3e7RnO7hP+NhSR4byfMwQ2UFDBZJ7PCHh2
2FdgCOvCoY6JbByMMZCfCNAsSV4omdntgukRRhL4jdMdnq2posVdKQN/tRYfUq1yhdhaldq7rU8+
Ws/2shtdtlF8OQkTDCADyqyfr9X6w2y0LtR7AA2xwInLvtqpiD/0rUK+SKYPzQ7mRS1ZkG5t74KG
i1mv7RnmS3YzXn8MkqkWK39vDtUBIeK3qSxQs78DTttqhxoLMZIJ+Zy/u1F+az6AUOflfu5OOC4z
i6xq0ofCVGKGOt4hCfYOpWNxr6zuutFX/13gEid81gdeQ5p9IT4j02vzEo+5YJISvSYe1atwsHVN
LZjivE/3ck2k1NVcNH0hRAPbDzJC7aWnF7QU0+adBfzN3VL9vVbjpl91baeiK6Ny2ObrbgGYaBmK
IA/puhSseG56FLVRq5oXaUxBaDaPa08hYKIgHIRIIyh7PnM1FyuFBR6yXanuOSQknYv2nZznMk+a
gWUx70oShht1pOsOa10d4v/Iuu6L4mqTQP3q2+W3ovE+yhpiEmE5waavYAwsPReVKDsUJjMaP4w6
IxfxJiGkbRCoPdwN/94T9rGG6qwSTwPyyuuRugbptYW5H3lxkU02WLouqQeqtlxm9ZXt94iSdJgH
a9+n4kWIqzz6q3HMcdX+ahUrHtHILlWr0YQ9XDlGUQMxGbBaF0BWHr3r2w4AYd6brEhKPx/tKME4
HwmBao0MTh/Nu8Bf5ZLXjF5v2ND2QTDQbq08LcYusHhkFSgvYHuVkaqDe0pcAtbhnmILr9obWrWw
7u2cFVt/8M0DdCcuXYfmbTi1zjc0RMJFJzaimMB9AEu9LJ3+L8JFkgVFMZHx+IUQ3d/ZDuDeyGJN
BTLRuNUvQVacwNdnJG3p474MVxTWyS58e83QNgV3PZ6nN36+clrs37hezqbTkSbAsWfD7K28Yxrf
jsyEd5sRircpTQThUWPC2gw3o1krcZHuQ0KNShpY44rd2cLGNI36EprncNVDmUja+WuTh2w43d4V
yU7PwkGaU+cfm3rKhJWWfzEIBY9qbJnnCswK3slvCFpR3o01ssbkIdCkCDP6ba0hQmllQF+qohST
v4dc9v0nrJWjdmkxCh0JXI/FaGWqJlV3kvrVnlqmxp3751hnQZsTgOIEnh3Iet03aCO8R02/jT7G
UiDySwsSLxhkWVSSU4pmVGHB4MGGl+m36XO7cc9V0iCO3nvH7drudtboeooyBBlUQmpfLbj/DjmK
wH4HqMhRYpXaJaDCB7uV+AUNiZGOlinZVAEeNUt5sfhxU7jo6UBGzvaaykR8cCuGidomRa7OSGUT
nBYdyq6WfiFCTq1j6P4nlj/sja/eMH6kensrMPDumDm6NfaD5zvIpmtxTOGcs6aAu++kT6whQ8oT
KmN6amrQI7pPnCpvWjBbPuTUfIqZ161NEN9fEwzP12H+t2eDmE2KQqfKS2kUoXAylTwR8dFGYVrR
jTpOWbfnycXQ5jBLdLFruUfiC54WPdTNoOc2z5BR3H3riQtbqLcuke6QtG75Xv7vP0v4MsAO9kyF
P73fJZbIMRXqbnW5QnjHaHqi7Q2WnvPW0qlgElS9OS0C+AQczuuJJRX4sGUB5FuBiDpad6GaNfgi
6qEXbETQ3Z74UcznvDe1exh3d4ubimDnkwwhCO1yBOoD+5rDUD1e4nTtO1UVNRzYCYF+iNXwwLAu
Xq91y15CvMib21mbcrsSohGILWsfFzqFX7xOo7eqOXD92VIxZEdHjCaFnI0fJDLhPN0I95oYaxMO
PNIH8xAWoWDy+gGs651po3TPhGbZR8SkRaUgrRawY0ES+hvfy1L6EloSNSD6wWEo7B3eklRKgIP8
96cSTGC6mFQ5my60QhLeYTLI61M7XjdFDqQRUCkBjYd1JtJ6jcZlaJPKV34yGBD89PKhDp1br+Bl
2OXS8KQj1tTzHALQXtBYzn8CjZfyeCkg/ryiUdi6Q+rLGuC7CEtGWNi1pVvINN9rxOmmjeDmsb9E
shw4xrItpc3UHfciwFH2L/1LUyX8hMH+7tjUBm94pLhW7yRk0s2t3/Z5TYm1vIuTkL8H1z5XQgfK
J8RbvMT42i5ZipgYpi2BoGg520BN767dNI35wVV9b86MZc4fmVZ/2CdFwWroLRzN8Jkjfos40yS0
rtTED/a4JBp6ZWsU8Y4QhqA+NfwkXlem1no/92NysxFC33BL7gZ++5gZr0QOgT9T/I0MTqXYbqEu
S8SayL1s7NzMere7sN6BqEcgPOJ/3+V5mYSZ+OwibQsQPgWkzVgsujFtHT0EBGs3j1FPGu/gWjt0
QaiLmVLe4cV3pmbuZTWl2Nm5YT3eGBoRhU6DNxSTs80pQilu31ibEVFu1oiUVe+M55WzH3wopooR
MJzAbvlOuiocD1Q55/KlE4V0b19+WOxdkzwQ0NWzMVt2HVKcsLk8Ub6L1zXvESP2vCyD8cSdZsZg
NSom4F4HvsvkyX7x9mvHQzqeyUwB6xfO2u64boHqEzeAVZYezrxWjDfsyhqY4EJK1bJDDq7C+jsx
H4/x43c4ghNJtuy1tb/KJbopnbUQduhF+/kfefW2mdqxaviGerMFX5LouvpvKtHujdGObgJBsm8P
33aQwedS1Qm9zRXjCHsiARZwsb57lYVnnfggpNH/l3ikeLrdzKFy/GWEpJmBHIuNN8O5HzSo6AE6
ZDmr+fFFLF2V4DYz6qyja3rPFAkvL65/pvkPXAoh8ECk7MJuPeKSuog40T8JkbtBXGeWfNT/CvaK
RJIL52jYYqriv3PhLfird3uW9aPoaGZNfmyFkcIohpqVpm/Py8IqUGqqm04GWcTT4Oq+gQhJWzmv
lUpiSO71i6W8m+OSJYiZJue2vgK3jGl3TdxIdNfhu1ARNxmHC7b4oGFb7iFFqP/m2xn5LyVaFl2C
I5ee4sFsXETBJkkgex6WmkoNrULrgM3L0/ekywbxx2vg8XLvZuIm4d3J0boVIfZPYNJPVqaIHseF
ZQndfcPvoIoXJnYevktpwb65EZCPGPKAZM48qlFO28xksi2S8SZMZ1RGNKXbZ/o2WlWFaApDi5K4
9B5vaGIOouDuHN82WsTo7ZNVFz3cDULLG4KjQoGoeC8QAkdkUZpGkKK/+qS5I8hetV62u7ERPENX
F+0PiCaLOjw3QWJs0aJtLXo/T4gqJeiptMXCeFKGEajZWqNHspRrH/LAgvmTHdDyE63FOUY8Tu4D
W9yqD5jYA//2bJd9HB30drZ/DkFVos14o7z0ov77bjc/EPwCZ4wXcI1SP9gRU/T4ia1XAV5ByleF
naz/6AsnHk9SemkiP/M4TS0x5JO6Pi6ydLOk49vz0MhmL/QtXm1wa7YjUiITO0lIgh0NFaRYWMXh
5ZSnJwqc7Mrw/QXVJEgn/MBcLVLMLy65DQ3+yWVYBCqIktlJgwpwTSnE9WaIbR9xhLFY3z2eVdr6
/G6i8qbWTOFssSDC0tdMKitFrz2EYSFodJxm26KUbTsd6FN9GVayIBjecZ+UCga93ZO8FBx0n7i6
IXTyvZMr/WvGO24Ohd2AdFvu6JBuyUUEA1fC8cQCYH49oAn3aNnAxgjnykdiz5fLMnPFHqbJ97u/
TL7Egws6we7obYV6XRuJGTvdyfn5oScd3Rmi+4HajMnlm5lW48h9OedQhuorbTk7A2gnYBCBHiV5
jw6FfkC3dFizt80jTh6vQM8/kUWf8EHdcgZH4TwnIDJA51TwOhKUgfJSxNFKwpSqiSKhnRqx3pnR
2x0KV2UxDIQxyuBh0Ix5lUO9sdqHDIXDRRUMqyKG2z207MACGMS4Dxbp1SjnxZEvqPyx7IehF8ev
d5pO5gAnjaiqyO31k8nM6D9HKgFvL+tsfEAYm1dmG1ln8Ij/Aba0FGLhB4e5fmrG9ri4UoqOvcq/
6BQ7U9NG46OY7iMKRYISBAxVpztvEAmKJnVSd5b/Atc28v09YjOb7QhARBN3kFv7Hzy9C3HIKrY8
KdMdgNHFC3cm/qFJ4MsfxwA8WSkg8vfsCbls2qrVI1thsKolpQvVuTkyBKEN20aiRwssa53bFBPQ
WlIsGxBJ21TDWMyesDuJA16InVyrCqKjwYhFpJx3yK0/eHY6HMGA/WtQIhKH/snZiqodzypkHKe7
2XUX3pKhtTqzY1Iym4q9z6gmrRL/T++UpwyzLwlZcppoOwVKfV8M4vE6iKOTwDOpK2VNMGGSW8qV
ZgiruxpdJz3ylGrN881Vh+ecHugldQ+GmH9nQ0qNocUHEBm9cy9GgbTEd95rse++gL9QzssHJ2ny
Rn5yo6Fymm4i9KHCRrvJ64+uyWWLLxP4MaEIdHkB10gkp/SfO9DbHrZtn59P2amrc7CeS7gkQOnZ
oSkp8k4ItBPWIQLweGeT/vFRKPOYBfRwJg/DqEwfwWYJQ+ah4Gvl+4eyW9n2UCMniVL+ephTHPmu
4sf7qnkfAqPBdaJTiv5H8q0JJUk8sWjNbbRy9YNws7xXp4siGT7MxsF0lEAGPDyDGGqff7tBCPFP
iSDvNC9XrUU/kpCjGNTSsfdp7ohlCNwbe1HZNLrjHRizBVBrDRolv6APpOLzo/eW5WfUgPqJJ+5e
vAVL9w+8Bo8E+5Hc3ue4mLAjAls+NXK1xP8kK0T+E8br5qBnCfgrYNf/lrsVnXA+SQ4n4N6gqX2X
VdAXPkxxPEtICEZ3DwNbN/hHayo6Zy8yD3aR5ulVp7Vx6PNWNfBRJm+VFAtYSCcLC5r+W9vJlX2P
oH59XTjXUsZhu5g08O+4HLFU2botFxTNG2Jh9S8C+l5LjPXra06nRhbhP8/nAwHAfX5zxnZC9rdH
4ObEdLjqGp5ytH5slR2ozf1MAO0+rUzJ4T4zHVCPtpP5O3XAs959c/zJto4HDNIoCMmQcOGDAimi
bwAHPqLfpM6TqyPuRHoZo3mVzm4dGln+8Tbn+cu9/ukzMWoP75yg8+SYpu4luTRSpQODIsmliV5f
uOPIWBvNl+5AvntQyhmhGjmPB+fSDcrlJ5+SUlp5uPt1wDcGMh3Oko9OIFW7F6DTEYbxmdvcCkEQ
iAJt10HO5SwPCRyGL5H7GPfF51D/Rd3eLTzVKwuakgk84s4wO9XzmUSiiOzQggZdqgLGXBqIX+Et
DSQhCYEZSC63adzRxFAt89wIXyAafcsWsnvx71CECCRqHFwr9rF6ECzfsaoBqv2M88wxtTt2Grm7
bY28bT3UNVhPiEJH0RiJG0p+uwK9b9pR0fQa5GWh37toNAxQi48ySTN25kQREGJ2qTxxbVUWx8r1
PsJ0NI4JrIWl8OXEphOZY83s3csiLbHn7SOixFtqMkEsTrar9C+Zd51CtuZWoBtJ/jjSQndYAVSs
ry1uoP/pmGAqz35c6bklvq0kx6OQBYniqL/8Uw3rRXlzrI/abAsC7FeRdwwmgs+Ljl4RYPZV8P1v
n4zB8TNBDvd3x8OMjXJGm9K+mqdXcHmT1Io4uqSmFEDD6kpSmNy2nch1s078arive9EW0BVMuevT
l/hV98vupnq+UwwTd9nPMbqdNcH9qSgu7qVzo0DjjLNCoaP5d643GSj3ypUiifgHE2E5BoJ2jUV9
JzKFCmsTo9SUJWbzsonB1TaYRUmtP0Q4SGNuutkTMCw9cgmz5DVI2/TZclaFosTyMuYGb+BvM7uz
3MSeAOwFgXfA0xMfiA2oe1awjtXb3Xc8QjOW7Zgn1yPy3H7Z55YNNj7GBycgN+5IP8qaq1kZJKii
JwHKahyQMz91wxAL86Wcht+ExzC3+QxVgNwFF1MkgWF9au1ICI5glrx62tESOeGcfuB2Yg5i3kPc
4VuQCCPI3Qf5fy2XKuxk2NeeCCwSNGgbCaABC5QBCEqV4cwzeWUBrggmCyF1a3BFn8CrxsuVKC+R
AgCW+6sz74La8ZcYeo321qz+D7N/8RAy4F3hM2kElXjujBgQEEJaqAKrQzQKZL14OlInMC31w+aV
M7uM2hQ21nZsPUQJIRwZ84lbMuNrT5Kdrmxhb6kcCZbDUIRvIcvtLpo7umWRn7QdXqhEY2tlbIKP
xSYcfcbya1zRKy4MLW5F2iKmA8usjrq2IHjmxgrHHCG5AHnOw9VJo10zJN5AwWH7ht034fVrXmqM
kDlD6YiPDZ2rPSeseSUpMjh0JZwHG5dXcmXja3PnfaTudRFO4JVMceYDCYHN8CeTJqCx02lIKYzb
4oy+142J7oVyEOCXVmbbIg4TKgqZF+WNsR+As0OpGSIOOkz5Pegt9f4UvAxRqvLsj4PgdiiZ5066
gffi6jazw+TSc+NclIrDMNO1h7yIdxhZOXaHQ4NsQG8GCdxIDJKGgv2gBT9PurBTlnpHX+k3JvPT
i9Gq+gwZiFSRx156FUgi8dg2ayN9a1UbDWWW8IhiIAe8tRFwHPaMmdfQNUQ3SCOXaLuiXi/iV+iz
CFVmajTAmgJSM9xYWmdEhZLgfuVv2Cyj7BSYVzSPEuLA64ziO97YXAYU31X/+kXFCFTfg0JAxrTo
3FCpEbHqn/uB0HnSimjH2b9J3qnZ214QOGgKRhV9vpEw+unUC5siPYMQjwSatpa+nPWNy6UCGN0J
maC/8vzF/fLiWSMfLSEU6XFwDc78QLmmPtStutOiRlO3d2rWFCYrQ6N2hWLspp7KCoq2V+rxXhfr
w+yKEFHxBTqucy8JBzOdjFinYxtz5Wxs0MuM0j6ymPdNpszVEMvgsr5T8XNHIia7TPMfr0pEZC3X
T2FEa1WqU8L6LVKJSIx1SFFf1Owa/tW7Uc0MgNlcaiw7t73JdFaLsGoxqjsTrvYkAAqFdJq1kORO
GfJ+kF7Q2WhgWR6oTMV2kYIW0YtSmK835qdCTJln0+JkZEn7ZRMlsPCdDD1SJcIAE04x0Sc5YUbP
p3hdutlIRi5zXxUxVHTKzG5MpgKdH5ksWI+Hbk3635qffDWRoZ54yl27QBMh4VK8oR0yFcwuSW0V
vkQ/CvhDBcstzeo+MS2peJf3ICnoJZ4IYPxCfiBOfYDplEvlrUQM9tOQ2+3gynUdAJoWBkBvTow5
hesnqD/e3BJnyJqAHSFYMYHg2Foi5aIJRQR9fdu7lDU/5gwlsT/1ceMnVBoDJLRA1qU4+ZumJRjJ
6Gj07TpNaFu0mg7pRuiBwdQlCrGHXbDY9OWzn5V/Pg5Rxcn1H8WluwKQi7P8x617lJ6MM1k1Jk8s
AxDTRHD/fMDZcNWlH41JCqAEpxpNND9zempMAFVTOCziCTZMZDbMKUhTU3/G4iqtEInzRfGjAqrG
+5S42ZDG4CdE+wh2DDXTFEWybG6rOlnLCHj7h8kRAYpV2Tck/NM+ysojRhr/vHll2NGFxafwIalw
imDQWFeyQ5DjPN6rkNinf0Jk+5LgZuQ6LfrBAx15bVNRB1PCs920TgsuMS4FJ+pscBXFZ5azjOM0
BhNFP5Vy6KH150UBDISS/8vBuxHBBJBuo3Z8BYGTAYYQB/QqDXM61PqOhqVqwoQYYCmfP1ocsjGh
dSgvI5zcV2AFGByGYZoE/B6eOlBFdV5qnLClc+zy0Qaeqfph3XRu2foKUsaZgJPNfrHHoffdrBdQ
SerU8euSH06HtuvHPFwwFAcK/Qsn2mQIXv5LXbo25CO0GRjoXfyJTKo66y067hccR6skrf94Q2Va
jrj9fZsZGi8aRBzBgMOHOHywIRKaTz2ksMBZGXe7/pgA/u9JTfvAkyqFdD2WABcP1mv3NL14WZn0
69HMfugKvIqQwDYVVpdm/ld6TlE05CeR6GUFg7JVAPFse4EfHSpfSrUbWEPD0LB/bQOGixUnLefV
e3SN9JmILS/sugjnct6DjVCH0/pezNzFJA42Vbwie9YbTl55gNF7gvgDzlZtchhDDsIjwM2aZ6BT
9Z9ZpxzsALG6CXzdKCSdo6L7/pNsuj1Un0q5/2YNYtCsc5/yinEVGY4Jd3LthKditoV34jgIf+TT
V3vlJztfbqki9MnYNXIXr9RcTMcw7592KUV+yTXkIe8jT9VEq/q+zB4NXzp8B/SZmrXwtmJ/jsnT
0Ah54937VKUXWg+7tUsU/xouyLL0JIyuB1Vh0htX2pLsY5gPhNj4r5bu7cAzW/fH8IaBA7d5nIth
6ORK+wPW6LgL9AOOipIQH10LAs2ogQWgK4SXt1D77/Zd+NVEFv9B2QPjsvvETpnxRRQz4emFYQi0
z3qzdcntb7O7+e0Hw5z/EYKHUdwCeL3B4bVR6lrH01J3rqEm3Q2tnMa774LGCpeP9z+317+yna6J
5U0Kltf50cY8tabr4rfzLTozAAXuYC2QyvLjf/kIf5A8chtb2YAmSElXaL2ms8caAw5PF/ZsSq7o
rkM2koeHvabKrLn3Zc6Dxmw6h6pWoofGhxIzwNK0mvmRMCP9Nn6vLaXLuhEsl0Lx93c6ga0GihKe
mArFepQ69n6Lvftl3QyWQK4oPMPcfqcPjncDfv5vKRWEz3RQv3jyP6bfG0JG5z412b8vxaU+gjvp
/9jiTfj/2dW//K0raASaCpS9244n9BmngIBbEYFTx4Egj1KSXFWBrUSkSZlyojqO5cW4RryvRbZu
SWmRIqZsP1dJKmvTb93bpaGpkt9Qbb1Jw2u2A2BxdkKhu3S/7/N4CU2Mt0m52z2s2eZQxrzgf9bd
gEutxk/hQWTMX31Zhrq9m4CkASCrHpfsV+59kkhtBpXdd6pZpzuNpFdYaFSzpzjIGhDBADtW9oyb
wK0tv+1kBsSjiNNU9RpvnftUkZSbwseckFNB/H9n/TcYHZTOcPopiKwi099QTJalDHO8NXPK79B9
hB7pW2oVK2pLQ9aREa9iShLSMjkMp6iIKWYkuQ3V22UUglyqrq+mgyPvIzQoEre7KNo5OIj+680F
HqnEAwdj21OFU+wpe1ckBYbAmkkaW/FhTWCeWvKyWBiRf1ttIDdVxwD7o7xIhj4b/TPHM6wbmizF
NtIheueGdQ0gn9hPC+/hlMciW0CSt/7N3TZoJ2j7Wek9bnInLCg8LVr49WoxmTcXqR8tSI+161WV
WEBG6x1KwjvZ2ge6Af/gQ+ImmCG7vbv3BVKC9GmFOmWqYxm/QUtskP2F05lARcJ+eiP2K1aH9DVv
CvSsO0FedcEL690xSu5JZgo5/TG3YzsEfobXaEVBDGtFKl3bicAbUZib3b94Jr6WdtBexkT57n7O
PFph5+id1JPJLAEqaaiNNGXCU8xRl8d++SKx90iGa+MPZy8EfJro18Q5rGXvOH11XxNjw1qUuvZT
Rt/yMGFNQeujSeK2Lvv2OUQkJYzKGVnydZ5u8wGkO6Qr25kkZVkLFAjI4OeDo212jlXFhEX1uBIA
nHYfasB9Th1LhXNeVidnfZFHs8NEPziO6iKMXhGZ6WbhEj085WTrxh3cUiV1/OsXiTPrK3vKeBZP
rFHpgLvE6J2gLI+pWp0TXNDv29ouYoLMeJ12JRgNln3m51sGVNlgo8yCIAyIfiRTK1cEV4VK/LN3
7KQ/IpmyA5rHw3gxVZtQcFSKEGeyZtt40qmxHyIR6O3P64+Rqbl+n/yV9LrRhKq4gaCMmphuadVV
CWxe05dhyfpWIgH8+/V2aMKv2JcjrHU/54egH6Ysod0gM+EQs1/jdAIWF8KPCqRQbZB1zxhNtjjT
OmXnBC8vX+oxFVejPqRFJiXotVoM92yPD8wFJgy5RcFgGXoKiVjXc1+j9Nn6Oq1kf7bSCatvVF8k
W50DUTOcBKzn1aeqnw3rAz4wk1wnVHCEZNgDVMtI4s4/Ey30n7643ianCfywiqzKAyiClh92hzvr
mNjZXH69bc0NGF5UWSfNFQ3cGu1KwmJMXed1ZcrWKPq3MYL9Knwnn72ssghPYucd8P/YIetvBBZG
ip5MrHnPP6t19BqM5eatD4xp0YvoYbX/6JiJfmlAK8xz6LogU3qZA46ebdxIL7FvsSh/b4NDMZgL
oR62BM3i3oM+WtX2KhLQlUAJptSPunayOF0dzct924rI+cTJiFOvu3b2OA4CkPWoYrNVcE9FkfSB
USEfGz6qWNnr959virMa0t3NT7FMaTwfC3MuHzQAlYZWRROWYWKg25wo4QsOqhBDCLHAg5qdHQqI
PhqBH5cumv26WQf/JeeQQpl/fp+bTfzkZw+3SoWKjyoP1gLC6q1Coha2pM3KwXKVfvsr9dA8hE2O
jN901rcDZr9deMqMyNIOWEd1qRHCnQZcsDDLG8xmaCBonNylvgYGjQMTe0zFr8ucP+uXJnxJbc7V
9UcEG5Vroh2xTSKs6fO3Y5YyihjnhCAMi5qUM9Vk3I+RZB98VCykzOlwWRHgg6yAdsy47CVRs2t1
MBbeb44aCi/+xqql83nkZNbLDtBqe2uyXMas+XuRhqV2f+QrhV0hwS8LTT03bPtfCJTsYp5vXbRJ
qJK3qvLkf9AGtBHb2+36i1B73D2ZIBGAakRK8yGn3sIwj5Z3e08lc8oS1rMbFPeRVGOHfoJMYyIQ
978Cj8xtv/p2S8r/W1VvXEq1573QQO3FLpCmR8PXu36k9a65V4XEdUCKZlWyNV2fjxYc+nrTmNNw
LdkApKPi34ijcjXBTXwVjQOFTfXkU/gnK1ckT3VZUAq80NyVYcYQZCIHAmwSNSZiO4uf67HkOivs
d+eUtQ8Bm9JgvpGmt0x7DTdQ0PxB++HMPULucuWOmFZa8J6YLNqdO7/r5zGYuSzTV6wRKBSK9nQl
pGQs+X0I5KTaJvG8aXnpayc2W19xif3TlikmT1Tyf3vzVbv2UChZHKcvMuwMmdr9HWjzjFTu1t1c
RDIU8dzo7qq2sXE3qt1TcWPZXRBUkDbvDhwn92O7MVTnctubzczRrj65puAXPJhrsbF8Cn3xtNuq
O1d11rfxogb5LCgUUkgdbs9kpfuVxE8j783wvk0LBawXTz+XiAuPIuaGknHtnKzl63iao9bkaJZF
fWnSuJI+eT/0w/Z1KuuFes0rP8TwUSu0oWVpVLq2AdsOtREOc/JsOd3iSVbgNLzG7GBeXTH9hKz4
uVKnry/2yNRYso5NAssLkl1DdgnZ+YUVo8d9eXSlJeWMyRsXZ7OXefyy/QUFfCdS1JLkywWzc8f4
795FZk+S8zJiFLFgv3m+PaZRiT+OTeShWw36i/u36+CTY8IB2zrLJgxDbiSpCVM/iumoCz3/1ljD
bY7m3162CWiXB280hUZa/NzxxASOhu9Kc74jOiEu5lx8P6gF+ni2s1z6t16gJc/H88HcJm5+Z1FI
ccbAbKoWVnkUDUYPVVIJIHiuJs/rOQ9DXPu40xKced+tw0ddYMaqQh98mBMAaOI0fpg0MSxvnZad
IQ78p5njgpWWm2WXoFqKNzDkbo2TlU5cCw1WdUBZB/DiGtHhAn2lCh8zG5HU4iotrr8c7QOu+Psp
Cpm95gJK5//xC4ZjvZwyeYNE60H7xCUKjYYSOGUG8J7lJX8GQiDd/2CQfywB4uNFJyW4kC56F0PV
dP1iyZ8skm50ePGJ3xaLvOfm+5neD50QpB/HfENCeRNbD+F/wvvFEJOt8qgZz0WLrQJZJ+Oe+98v
ewU4033JD50yjk6zvttrEm4dcAtQGQEQcPBjVbXie+djqKz5mANa8KmUku1dYdsKyumTNlZA0VD7
ds82IA2aHkLvM1GoUvGj9ksJ2RY0tmDH95jr9I2ACqvOeb5DPVielfvZ6Dj/fTLVRDD0JPTJ3Cl9
k9BqWzrP6CrijqFL2OVMpSLOp99KzT2kvivqvBbq65jcBrb9M30msggamEnj2NBSe6vXbcXGOlNI
N5xqgquxhK2zxMLQVTu/ZoIhlfTkYLtnoYueLw9MqspowhnXXecah5vcxgTxOxHO7PklLqh23UXN
y5VGlOTOhQuzpIpGjJflgYnE1/B7esflcuYMp4tOid4j/f8Hm5LPP9ZR637PM1PpgpO/r61tmria
/pAHUlvCfNtEVb8rHHG+5llrJ2Ivrm6GQM+MHmDog924P3VW98XaNH2EVeQNBD8ODcKCiOq229vp
MjNUfNo/mr4N9aXWO/QRs/90+xnay8TcPejVjBkuHGGLYHGziFCw5j/0e8nQZb/3Jgg7W2dkksVU
sTOM8BUUe1Ohy3MHrXiwjYsLJIjXmhlYkvRh6+MgbG84H5wlvt0O8HzsVSfTi92evRdSx2OKBb09
wzyr13IvTUOpdglcCgVLprSH/o+wLjyHA7q4fBm50REDaY/0gYzYoKeNV6RdwZ9K7VAYV1y1ys/8
1ARf77kJiEj1H533Xf2dY1rtxfjpYn99ozZXc9OpMibbFChFl8eAtL8S+K7CJPP01Q1KpjFQ7Z7A
72yaYrdQEYfWnS+4840ETwxGKE3xd57UV6U+0sDmC9CXL5RSkXXYhxrQ/1z1PcmmeVJTmni1HVop
bWtnoASr0vea86XAscU+YlDrRn+FzEgZnLs7And+0Nj/ROK5vHrI/Kn31/CV/UfSRG+Y8LiqUJ59
w/6FiwQR1cI5XuO27wmz6UONpVWmSMzi9FUd2+fKrSgO4Or+l69L0tPeGXLHe2c2d9btTJAosmds
/D8DDKw0aHtP2KtEBlJOaMBD3hB7kRqD5Tdxgr5i50yft4VJoPKhV3CktP9PKU1ZU/uMRQ4+o7Bt
x/JCCJO9L7NQ34lOx84eSKICQ7eoNAgP8XgPNxKWepp0zEjvi+a1knnxlmBrbF1H/cMere8T0gFD
NOv8sMOz6K2ldLQqZNRGmjsFTmuExHJfPjbcYPOA84S1i2DjUThMldiPZmM2UsGM8L1mUdwnQ2Vh
CYFaOSJZXvxROLyWASv80aVUsE5Q+SSIy8zLdz4QLS8S3pH4//t22iPw7JLwCg+Ya4CNbCGohcWr
ruhbeVdAMcgBEP1KKtc9XKGSlMOuQngwko+qbMMTWYG57o6J4jFrEm0VOv3cmOvTMBSIh7b7Fgdv
HvO8/CkMUE4gfRlYlqBU9hbhuhK07ju+Rf3a6j+U0owjiHvPau/82MFr0FlJ5RsHDh68248ZdxH8
4BTn2yipbBV+KRfm+e9i7umd3n0Wa+T1VPDG62NewZDFm/R7guns0i/r0oRlHqCFF7I5nofkFqU5
Jwm6+YWDD6l6VYnhYOK1DzrZeOBLPPHDwaNVrIYkBg2Fgnjmxt6ysP9rOiLDD0TzCXHxyBbAgbmA
0qubrEiLETawWYW4ejpRSULLEDopphznojOjj0mI+hPd7XURlC3M8QNIpco6LEqQVK4HHqI2iA/8
niajJ+/3NKkLvF+N1XTNnsCNh2PHjkAUX+nozov87GwxTbTM5bbPwXgqjK7bWVWnBOqLRf8r3OyR
IAL//20mBDHVQo/QFYOAuFCLeDRX7p04fLfJUzJyzqHxFUNkEhT5fSFX6xRACZcvkcKx3Z3HmFJd
/IG5nWclPao/hmfFsu2oko+ZljNeS2Dex3qttnKDlw63UthEDAzr3z/FP2JH1q+9j63c2whZjsRZ
5RpK3mkQYTNjKIxK89ssn5zG7+q4JpNkYtOwv8aHN3uj1Xu62onOVZw+p9tkYGfway+0Dn/MqLs/
SI6TZ5zS8VKgM+Y4PrTC0iQSq9QEz3/Cfv1EGfpaKglRhZkEAbBf2UCCjVGWb4Uk+S5syeqCMuYL
V/SkltPCJ2M577WjWyc5yelW1UQffMwGFG9dOzD/JGp9Nu0BaVguCPGJjZ2+9pJpEEs8rpMotD6p
hXrVAmzgtuCmoFCyuQcGnRVTLlzhYRkq6MkOfKR1ijpgRWvfhxOQwEjHqfK0DFx6Z2RH7ASCraHg
JDd0/TzCURuZYbO5bGyUNpPQbLL6Ye6KDWFr2V3dMmJiFSQOyp9Ih1yr8r5PyDRGWpwDgjkw9AkB
ceX4z5HevvMdeJoz5YvTwE7eemxFf5Pc8VdG8DRz2lI7b7dOcqkPapwagalFVaFnh8HJ5myLyI9p
5VaSRjpGefLww4to0WYd+48AOWRD+ZIrIWmvRZhp7N09C7PSuol/nGoMBXlv7HDXSBMDHdB/m+Lm
BhV+f6FQ2HlADkuA+jW+5F/F7YoxplabMDeGkCzE0VdCgEXcvHGrSh4LkBFvPFI1ZTf6oi4nNDME
26P3utOKrr5ARqcDjacXZAs5HImpR9qgumGOz9DsQjC9Q90axWxtP5oPz6d+E7CSF35TQJOJScwr
a5eVJA+udRl88QkcMf5CVkTDEF1t3bzD+bhxcJ6aCJX/rCjxk9KW7VA21NyEN/SLl4fM8CBjl14K
/RDNvPykP7odNPI8wUGNi8eeKN+LPBPnbgYdnZeUjIn2XF5KMYprpwFTNAGhb/953h7KomW8pwn8
N8v/IEci5bsNyfeGRV8R+xucsCZvabI7eiOWjtMh0bwDshu46i79LUyGwGgm3iLPo90FpyjbvVma
wW97dchT+wnbJGSQSEhGqI8PMh4HLQXgkzWD64XGVFGZC89sSn9onmXugBKTHT+ncWyRKMYAdJE3
BPslwwUagZ2VKZY6q5RacZQipj7E+E5RnQDSuk779JE4mrQMHFjTxqir1W+4fdJv5vB0d9Y2cnrz
6qtLCtkSc4dWqstsRZJjDawA4rwLAvxEcUY4BoLfKjxQuHPWGLCngAxBy7t0Jto1dhFcgYCt6yyn
c0kcAiNjRPCOX4VayDPMX/kVlZr8T8/MAZJBB1rVvrOEWAZPKmSyFnrz+epejhpvXCuYi2ljfmD9
MaAcLVnEtta+P+flrUgzcRzr069syXCvCyKxZLAvv9lPDvqSVIYEGD4RiTIDqhhfi8wLoABbdNfh
2zjICOfToS4BEArY4iyMNhWgyb2MBszTdIZALZak6Cqjkf+n8DoB94Vmf7cqgY8YMc4cDavdKHlU
LEzpDg449NfxXpPb8Ee+XrJ315G0ae7mfuSYz6nMj8QO5iSLjvBXT+Vh4CJTjWonGe2kyuE3jczD
fk3nyK8jGLF42fwJ+9l9bATcDOIABwQ27tJ1j3WOU4VN7nbDUch3+iQS6s8ujDDmdX0PsyV+/qM7
5LReB98BjHYUqskdKzKZ7ydPyh/CB1yK7CwDuqZi0XBfg66GMyYW1Q8kELX/sWHr6kjCZchiqYQ6
CL/Vs3P5hJPxfWiJHs9LxoQE9u+UFp7S3oyg/ly/xmRqN+jhTsaYeqQO4TX4VCuBXbMhmJ1T2N5Y
QSf5DmnCj1O/nuDKHAJIin92abdWcQGQ2gFafm+4eK3quL0Z0CC+Az3r2p0yCBaetci1otQTFYVX
Wf4XVe2p44HyxegxzaU6hsQ/cT74JGBQfPeKzfM3wZyuVm49mJ/86S0tOT54ChP+Sm46dfXVbs1z
prFQ+Dn4sJg9dm7RmxCRh2bspbN5x759c6xqy7qnwSMGFFlDWMhvIRQ2Td7Wlogn0XRrheFUMN/A
bZ+7Eq2+nNVj2lYUjQNSB97wn4g8Jk+qXyD3BM6MOZbftytCxvhrXjVD9ppWeWSia2gJ82XsMa3f
zx2HQxFZKs4Eo7+k0923kdh6UaKclwelFpLXt0/cBrbqmsulFY/9JIY2ujrMMce6PztgLP+TK1h2
IFY3geSeL3JsEjt6Thd5l/NEJEaDkp9W24tuo7t67uH+fTCyguwI3pVHML9vmhj83OgR0weO97L4
/0VFHKG+WlVq4DOXgTC0QjGujCRZTbj3kYpHZZEQy38l26ZDF5KaVlIBVu2IylseUWO5x0C9r0Fs
sNKyk3gyOamjIl6sVc3x0GzP2lLRVgLf5VsLu7DzjpYXNt9nW+HFO9jCUc83gh+SPyUN/r0AufiS
eOGlgyrXDBhnn77gcLyT0WPp+rTmbuAJ4NNVvG+DW60goekjHclJ9L3k33nMqvBidDGmKOnXDEoK
DbRNOYlDyZa8XdnYG84QsuEyLLD7ikY1s8TtsKoD1NO/Rh0dSCB3aZT1SbzSOYuDiGBRPlvi6yJg
/OkbOkrJLl2uaZq85zgdPDMlbd2aX6LZJ/M8kumgLb5zHwaGwaBx1xjSww/tFe2iparytcpGN3Kd
eeGLwrmVOTQUb/LIasZa3UkDKny4IIs1PDK7Qxd74wmD0HZgjslEkJXAVetDxo8JnM/309/u3IkL
0fc4oBvI2xKidYTjhaV8udFEwYLj7W3UWZB31ttX5ne+c7mnk3X1wtOHfu1bQUbrbeewaTv8sfEx
lrP8QHjgs5zMD7VRnRXGDnl4zUnHRBWT5N2bSBKcoydvvN0CeaMPGA7kzI2ygPEfW6pPryeKsZtM
vjOCYtECtSDq5/8oqCdCuASR2+tn6qMQ7igEjB5L0PWb/cbPfgVwZkFDCsS+kbO9NxTBDk4FnKM8
Q+V0U5M11Rlhi5k1dgFlGulpBiAO8EiNOuoGJ+MEoO3J6DoKjAwUKsbo6GwlaL8rCNgxMibkjDRg
I9ylzm1skV4QCadGJ7gCpuqje+yEQ3jT8L4ITjMKuE2hU3iZhf/t0yFx1rDHRb/yfeTHrZqxHwK+
AoMFQ++w/cWXwNR5i2JeTwB1ZHdUKcHIi1Ez7MTlIfAE9XNdLwY7lNiF3xmqr6wAc24DyqJgzDjd
JPdzan98gRKUSq3IqE91sCAH+InoeJgvkBQzJbH+DQ31FRn5Rx7Q28YZrQjlyjBhLj5P8uqeHzHN
7FzIbs2zwcCimsva0hrGr49TNFpNQpNg9gcTdDyzPDnk2PsYqiiAhQqITW1a+hRA8a/Y8t9Nc4xb
tduZ8aK03Ua168CI+p0uZH1rzRJ/i0PaYN4rjxi3GrmPJCP5iMShJGBd2CJEKvt6oOwbQWet1WNC
YpeP8Dw5HcCCprntoHmfkWOKumhYylMVDTkZpJwq4aFOb7OsbWrwQGlsgSEmzj/qGHeDrIPM6APG
kSMw8tAVy5FykS94zZgxclFZ8JH+GjXzCYGuOdz4Y0hAksbmKRMWL8Ypa4BAdpC23PRbgwrsA/rD
h57dREckFT1KOv2EXFwmvIsXmURaSgg0ps2KlBQjHAXAdqtwVHZwleJ9iskTDpT/kbEDhMS20HuN
rhoxOtXqKomyPOgoThxVp9Gh+NlJHKpyqtPLGobL6vBYNR+iV/7ufx7XKbGLhKq7DCYq77fv+EgD
6KgMOq0bCKaNqg666O52S1eKZUg5jmWmKBXQYgQmC1Dm5LCOktkLmTvhOoFLUDAIEVV/OIRdT+3J
KlS4xaES5w4/MRB2N9rgzNT7Y5K6lrjGUOq/LmjDMuqNBI6uxlOI4StodZGTdoLZxo8KN7zxT2Kx
t22MkFI38cXYWqnQrDl5Lq7oVCQyVbqADVq1oBGrswrYO7ZL/q6Fh2D2OeVDOGihfC+SWgmKEsIz
9K+2LY4OaQhSioWwdjxWOSpSkFeb3cd9oYm6lZl81w0HntEAb+lUlho3Fbj/dSZTqakDM5lY4f9t
qUb+WQl4kBH9wx+DC7inCKcvoq5YRc1wKQ3GMWAVAStYBUGFG9Bta2F8lhBXLMa/ty2KM9R2Ns1d
zA2JCMzgauTYczZ+sZPYhAHg7cxANjAV3FWNdlERjrR7To7qATEVR7Jg1lOcdFnttwsUkW1ABn9P
vKbkBc8tpp8Zcgq6wNqrfnw03XuQzjI2SoxaTzg/ro7YWdP5h1PffNPOFC5s9YbJlwyt+/UIYDzO
JVU/eauXNcPochTTB9RuV+7/wkqIKYQiuzlh5ep+Z/FpRm5uDMWYRoMP3OsEGERB2CugSN6XhG1U
rhrdkkXKlpZWOyX2FOwA569bu4OczhcmcoKLpdPUXoXjl/3zf1+vlHf1facTX6Xpz3CU60E/GT71
Z42yBvc504PrXXbT0RTaf3tQDSH4j6xRK5kpdJY29OEesfvoDsZTNsuQcQlttjrDTQqjW4Qe/xaD
nnWoV3lQe9efxetZbk4XHnaPm0zRHX5oJrxVDvgYiVnRGH6pauo4fV2m+vEkVgYk671WdR66zW8U
fQDqvEt/SlDg+zPGF+v0/p7HfnpF/a9wZZg0ucTge1jpcD7nGJxoYAGhEkg+vQ/yfofkTaWs3K+q
tIMzKxz8ruGSQt6UOMwHVbSojpMMLqrNSNK79XR0BPc84ZnMn+LTcYgsJwNzBVw2vyivfyZa8tBU
YWxLY2uitZFMJOZSUdJwm+8fx0kXQGCDvxDpGfxL8muBd8sucPyi8/YRMrlEr4xglWwMZcVoZdh0
5n3fYrlEO2Bu0rsvosnHOSF1j0DNBkZrQBbjVL0r6POBtjdPOPaaCVFVlkeAnEt8hcOQk1eqG4kT
MP+6N8FTm2zldKOkXLBKu6C2cP7qf3v4nvSm3GyS8AW58ouqmcY5db0K3aSnUEMtbp/+Z6FWV9xH
yUyfV+Ka9EfPFcojDZ/ncZmE1qJVcsJtjX9JFnwCKMBZir92YPCj+WNQpRheZLgYNE7WLGy8KIul
+/8/rzNFNN/cAGh3//+QYsROXG0RMrIzGtqgH3A5GdHTXxJ2vLLlCnSMN8u5aLAJTNeAEf36RnyY
j87luFBLWRJnvomFtE1FfRBrnpVOdlcZdDbptShrHHXGsR2GcRFTh88prVHDMZ8qSqPiY61UoNwp
N18Xi/iT1nx6eCvTL4TXfTdQZywoCp6GjybMC7up3WuOQ4lNG+KyOrQ2vAsNpr7KFbNGi8Eb91I2
cBLI1paredyXd3mBPqFlPKRkXRDUZhXQQ8rDzXMq9OUHzN3QUSlDjX0OwaEcA4Zu5uR4/yHmzua2
hajdThSjypcenzbpiB7Uwh7CGxH4a7/0B2FA+jBo+BcFzyCnzpYRmMVx07UQV5UAHddfh6wnqBjV
uir9eZwgda0qG7mpYoglRCk7gXQyKkh+f/z3BD85/T+0Gs/OMPwrt1llsXRYmlkHL7Te76+iwOLI
l3vAvoo7p4MvB6dvyhgJoAIcqJG05FgLhk4ClwXXHPDHwVwPVHsYhb7CBFrqP8mJh1ynynW7cQnH
2UknMNZ0rhbkzgHWvYbRhLtLt4JaXhvZbZhc05gM8BKUxbe6K9rzcpgH/xK1Cldi6OXQk13siAPQ
LyMsnLc5DUcadeLs4ZZG/rwvG+6jDhSp2oV7HR/t8OQ14+h2pl/0nkRuPxKZMTA0XRMiCruqZAby
9y5n/JT0x/ho2pC/cdM3o1AiSlUwzRAX30Kdz4k9mudo1gouPGPF3t91Nlc6FSIkPpePD6H4eLC+
s+/g2KmH97shpdF6HSy549fkvA6KsTZnH/2XD862G9r2IugIjQQFyAJSWInzsMwUD1Nq07A3jdr5
ozQxb6/G4+Yi/DZnAxa3adI4twvECGvlccg/73FBn92ESmhvqTc4ZxIfuFsT8IM+1e9wqVRIE6iW
YmCjIK7UP+pa4Z1FJXCF7eptq9tvq6vjl5yLFuAVhFQkZRHr2GN7IJjPzBxiY12KKfePxaLG8H3j
0EeZWlpAmL1xEYr6NM2BJd04M/zUKkcpO0ol6UkxkuiucCQRy6ngNoXKEhwBfHx+BFxDtYQNw4Z8
gO8ADmh7pLjbRdesvI6A5pFyw0vjGuGQwGoCIqBbwBzsNqzbXqT+Q+JSmauiEr1HDnkzaQRk16ev
6mMNht7zTi7GCJOCdl+wH58/2ZTqBhfBgqf+Hp2p1KrGvN+kqD6mpzndt39dOW5gfvlz/v/Um/CR
CQK33C2D9hfpQ+MlXB8I0vn+OHczqOx9AQI7rLwtqG/FK5pQSV35HiQK8hbYFj9iLgt8gP9A6huq
HOxbMVr2sFfu7LXuY2/wArAMS53nKOIwdp6B9DLc6gx6cUXO3wQ7y9hrpJh5SoYcFwKVBO1rtuvY
8mncRHT0femmHvUZS8jUURKBwKG9luuV/O8sXdZGVlPkAO52nP49Q+QRfoNsQZzqtFgJ2+22XNha
G9bGiDaSRapMcGavNF3TFfMq2lv2AK5dYflO6Ek+OUE+D6gplO8DIPfRAgklEH7W6Eh19MwLFcCf
6dj4Mx1S5mRN/cqIuw+TCltSvXq7mxIKKA64MexIPGEGXAjP19tmiBN9zuGNqP0ReCVavuGqGNLS
Pyy+yKhnDfv6X6Xs3VqZKvyxTsMUJFV01mj2t223H75JPhm1u24yG6kew9tnYlRechqxzXG7sg5R
d5j6hBs8f09/6yhZF/JfYdVVbSdkuCPlHSnNocPTWhUiJNsm4QH3sfJdmlzU/bCR00Jr6tMgNkpr
0KvueNglO+AB0gpsrG6NvhTZKYqgoUPG8TV0ooxnzdM7tSwQA7YVsxU170n+DC88bOMb4z5XNPPw
79Geqy9dZerLtT9Uzb72zrio1buTbO7jPGusGO4R6gBAamT/VGP3WPVM3vO+GY7yU1caxm1n2Vni
mBQVKh26s8/MIKfo3llXUmAAiPVS15hLqig212fXLAIhfQR5FVptINB8XCvAmdZw8qPZwU9MkhtN
Q6xF911sIlPP/1uzNMc3GJvI6HGi/2qrLYaN5PqD+p3wpabmpsQaotPA8pdK/nR12XVUkFRl83N7
grOXX0EyGkNz93joXnx6UwRzrviMty8O+ZXAIMquZl/tUfLCCDcvcKS9yjQu/S92XGxW+gu2Rqqk
w1/6tVcOWVbJFgMG4GAMAAmrmBPTPwd0Trce71en8ljgHH/mDuvhnutOAV6Sl2rHNoqcetnGdlwQ
7n4rvnQgmFppnrn+q0q2DtJP5p0yLe32VIfWOLiLvhaBZHKgiyzo+EM9/3hyAUzMC+RjgQKk/a13
18Gyi25HtdpM2DHwtooWR5PUD1rpjtbsL62+FbmEsWwv55kRk/IT5/FJ+Fm2iqpHlJUKXvzskNl2
+Mb9yd//eEd9bZZo4s2dHDLYcLUhzxOhqAVKHhQF8UA1pwwY8xtS/DgKcoSiS0/VjGfBBiT4rU4O
wBKIPZTnKxf15FyIHkpzCzgqxqGl7GcqeHUWmcpHAR1GDNItvA8exA+cEPcbpQYpx1EsWse8Z7RG
7nWizKJjvBiVCBO/z7MhQL/+jweb7V8gt9J8W9LQ6yvpi/fiKbUm03xTJR/q+55MBPFYyquXxi/B
QL9LtMJ5+wZXkEC4DiyRfw0S7jbwZNHsIeFx5vhXVxupRVBHG013u7E9Jhp5q1O4vEQX4JUnCeai
avxxJ5+u6xzFBjxVp/V6BLuuCTFJZAVvAKYwTsxcvmxjUmzJByGCnl6AnFbo4oYMJuoXOZE0dTgO
8SQleMABVN3ApIYgHW8KJJ6o33hrjA6/uZMaiZjKXB1XyEobeY/0MY6dCrIsPhJYhBSIc0zkWFIy
yb2iRpHPdolk8h/vgaLWGV47Z0OHnNCDZ7mkAYGLQlmmVim8UrgiQnrH8hk04khlFEobSanXSzw6
jpm0PPhB5xdBJ+OQkFtgYiJJfC/hIgw9F+0f1speO66zG0HQfnZG0JrI8Pspt8PyEF/+/8P6EvEL
hIHvJrepEbO1tmIDmPWLvqdWvu+N9IGfiji2pUn/nsbp+SZPlOg7An7jxe+LmTsSRi1jsZUbPDOQ
enpz4YQLHE0jSgd/blSj0NlBNbZO98dBk11f3AajdKuqV28lesDNpchWtSTZclJ7OoItIhyGIwW0
2iJH50i0UthR9y5JThRrWTVz6++lHeUFfrSWGsL2J8r+uw72Z6okUNh9/99O/cBR33SmJAt85W/j
3tM1qN+MRxOv3rK+OAGYPLf1dVdNH6H4UH3kbgh4W4RNwvn+Z+pP9nSw4Nyyv9BduVKFmdjODT+w
dwyrrvGoHpmnhIM/WWpT/9L6jDJuAjo4RErtnQ0f1rIk2bGEvYlrBrCGSzComwey8hfOo4NCTWWf
wAloQh1pLI4U+ybfAEXAT3mVmSBGZe8qEa6aSXcwwCnwirV1A8ab0VX0ye0rjZ8rEHMrobObsi3T
pGBdfLxPsfg4VqhS8ZX/avskyLbz1X5ZuyctF+XjBX6Meq40RB0bf8k3mX5BGFz10hXeakYTVvh5
PSDvGFobhlGTdAzEw5AZoSx+Q53yVOZENjLFXxuWvum+nYIFyapXlj6QnSu+SfycUrx+8pBwnOya
UwVp2lNjNNgZ9jrVS9JZVw36/mRT3eDk6QAN+FXSVMrKLGDFnntcJFiu78CoADkI/SH791T/VcVD
oyVGT65CBF9RSP4KLicsu+7ByriF8ZvVlUNWRkzYJV6jCl7iSYfAZXm51j6JpeBlUCxnlhjNwBbe
E6SxkI1K6KtqGZ7788o707pM+W4730Tm6cp0BEMcQF/zTy9vtFfSlGtMOAvQ01BwthZPDIdElKvy
oNqCuDYDFhb5dvf67IJNBepFEiJLtch8GknapYFN6DQEUUp39QJpA4Azcblbs5ICWsRFBJVmGU81
4AyGUE16aYOUp8q+NjNuIECOTVl2HLU1mhyGj6lL389UTWQ2Cxthl5RH6Zson2vXUt7MzD8Yqowj
pWIyo+RsYGNt8e+eSVpRV6XVDOaQ6fk/EAifK8H0lE/3nAvXizI8+LWfCSRwiCKUKoM2N67jFlUk
CcwGaLJ/8DZdNmMc9gv/qsnG+Y3Fk6yjcgTHrlasfB2lH9Huh9snOpIbgbWcnwJ4ARxA0HWcKWXi
Ex3CuC15oRm+NOd5SeTFqa31fQ9GrZ1tlzdeAbHD0BtLPJbSu9ZHrsgDAJ2UPff4TtnNXUkgIsui
9apfHQTxgyeg8fw6HwifA3F01S7l5fW3QARt8ZdbhUJcf15JkvAbFxihZXxoFFAhqA2CcHxqXicr
I8qIldkrtWntHOSliBW5YVZweuj1GdG76KgZcxCDobZ7K3SMYdtFQc7TWxpb5dlZ3QZBtXrMMfdA
vRcxbnAwGBw5yAF25p6Z9ZiJLZUenh07y6Lu8cuSCGI6qA+xMxpgy/BE7EmbVowxSgQpuUliAU97
QpTle6h2dytKPIIzCeaob4jtL50NwXDmC8+DMbmPfZE2vn17mdJ219e1NG5CKUS9/9UqaXmZVony
Bn1BWtPZqYD+ptv9Rg8NvmvB0U+YWyLp188pPFfvN25z4FL8/G+TgSM+z49UCaLcGS3jr+MIHpdr
D6V2t6KJ0pKQo4I0fnf6JNSrs4HDpQ2O6G+8l8JCAmaCK+f/V8L7JQJIJaCOlZ0ZnQkXZ72fJbD9
gB0UHAcDWvNutEOV2Cp34Nh9CLN9jygZ2c90iKPCp3GHPWztM3LIWYpH1AgfUCRAIYEU9QiE5VI1
Ka1BQatrfGBpMiIuDpYRTubE0P/k0Qh86fYzyTZQf/Hh3ZNGwyYFMgCrfpiePfFKOIRe6uHjDpPo
d6MLmZ6dAiDbWU2fl/qvM7mswHh/MpGa8e8Xj84PzmU+uP4P2N9TFmIoYzwszvAWjFYJFmBB+OQ2
+hlz/5fHB26EN9oSgI1vxzj2RZzG8WKk3SqFBjaHcxOTOWLwD2b30IMvapTOYqjVLbNYBwLEXQc1
APFIvhO1OP/CTuDNwBf+v6vLu1wewn+34W/G5MEnSRCaY0KmaOSoyiZjt7ZfX01AbZ3hB/iL23gW
RSqopXSWmHjEvQW9aVU9ktmUVc2yA9i+pY+symW3lrVk0BCXzpNDe6aeyYpdzAkz15Xj5dcGboW3
llttslvP4zY3VM40oO6/3fFDzxF8ezDK6RnyWQd0/N+pBCLGi7w9dboz4zjU9f90DVKETsbnV81K
w1hAIp4JG7KF4GmJmIxKvJDJMYbX0qNGWWHspqTGFD45QWRQQMkSvjXqXSordUTAbccg6taeh+j0
kOsYcEpN6Za9Q8DoRpnOxkfGw5LSm+frhy+2FTe+eWuvnqvX93hovGoePZGuvH7ubLK1zx2d3i1d
C0Mr2D0Latf4bALHVMWTYP9EllmOvJsImzUf0jv7ityl91Xei+H3Qcu84R84V4bLHgfrtS4nvYc/
98bQzXDH9FvIc2Nm2PiWW+oA7d/LrjUStEe5ARAdDfhRkUwArUSWbIjzJQjJGA8K/+XHEUyrle+k
d8MWrKT5GSb38NDOilj3cbbIzBpZZXEbO86cD/a8aG8HCMgMZrg5Go6hsFetAaOfXIMELZyAH04J
6Nb+N+lU8vXkrc3cD4y952xv2Dz9+yTCiqajxmkEALb3pZGtsfNVc1pB9dnCA9FWrA0xIWLNyMig
5xQRw4atGaSxJivNq+msG7TbZmHhgfr9J1SQneXyvIppRwdLIMwuVbhG5qtzLI1zb1GNGY51yZ2t
lvicGp40CGNJqpSkzZkeS0AixPEPYRY3BlMb2CXxtG0X12baUXXpuA8TGrpNx0eziremoT8PchQG
VkXF67o/hWwTCLa+PxaLLUwbXxJ1DH42JT08MSIViNMsZR7I3wlclU9Rqd8LVLSThd3BjPmnwKFQ
fUBGsLC7zFm5gDAOqrC3EYGYAnaUt8g3kcAkJL2WZhR6jCjSIEowB9UpLanFYcOpKMwRHnRrv3T5
cLTAK/aVVBPLth1rnuINPFMJmJT59eMkmwnw8Twk4SUTU/H7FRT2FCD9nCQR4H5kWFmFBh2PveWu
rcKRbAB4NbucT+rVNMvycDMhlc6L+37bRglGung9j4Td9wUmMc44Z4045N/owUYCPbkumbv/WM6J
Dy9Lk0081Ng/wQ94O/yHJbZH9UfkubZ6V48LSGjuzfy0oMlxSjP353YQtCv9EXMLM/g8xTz/kcmw
tKIEl7Qe4dvin6+IowMgBXtKERG773CHnqenHoRs2Dyws8oK8Y5AKBPkTxWaKhYB6Xz/Y0huOURi
+JymLWS6kDqXrzazBCyFKD9yZ1+4RZp+Hl1HSIY49lq8ZUDzDQ+KV1MON2fg/9R1GY7gcHh8QjEq
vnJyWHq+vLOghB9qVTUMfDeWN/P6pSfLq9WkkfTmusOtMNrSx5C8Y7HxPOJb6WT/69DZF/UEWv4e
aWbtIyF+DPhEvn7Zh93x+pnm31n73tgCfd5IB9Q7tvwtNPogCcAjnf9VaTdvRJSA14Ir+npfuL8g
uiYTtw3ADTORPUxlOuNilR6C6O0UP8aYP9r93TB9JLdwt4SO0/9ahUn3iJkY53e/auELv5FUNUdn
Qq5aROGFJAqaoFGQFDSLGHEdWZpbpuzdjnl8G7SkwF7qPA4Hd1tBlJOB6y7Wm1Z/8cmYWtdCxIyx
Y9z++5+b6iww+0KnJhv9twhlCc9Oesl4yzq9olMGXi6UxRnjHJJcNhFLtQwCxRmGP3lNpximNHwX
C/KNcosqfbJe9DIrykD62xi8AeuGUAa+IsWlt0VVArNJpRGAKL2Sm38OL59whkbm3M5Qm0mLwSrb
r3MZlJHcQQaW8JOtxWzjjLLVmMtS7PQag0hqxLQxLJauUCccxW6f8G/sVMGrd6B+0GMPeh5hJiW4
oWLPSi//EPDIBP42EMsq1CT9E9ANfguO2FfpqYbSOoPi7fXZRRaPq3uj8tjE2fDtrdUoFKxtUkR5
WLtPwa25DK7HE+6PgwqV3T2iWSPQ0EIsJU+IZm8c5DHX0OVLkSoSetcZhWt6F+w5QebEj4lKXpgn
V/X3GmBT3ovj1oMoq/LCQ6Ki//j5wKXYV69HDcQ8sozAhzMlqeTdhYplLZ1aN8D8Z9v9bEpD+2pL
ukJ57Lw6q+nk/yNgbCaAe6tNSqvIGPc33cfxhYJ8RnBKmhegBUFbbGOjcKsG8EO50j3McI1Sda7b
qvkQ4UMYPk9YbRybltEQnoWr4MJJKEYQRyL7YO+UFh9hiVOy9deVOrugWn7HFuoQz2baWnlfWiHB
QQMJoT4ftpS7+LO1RH5RL8k210gu33Ko4nxYEfrLxONrUF+KXfGIc0WhgsE66izS3KBX+/eGW5df
yPuMT3Izcs2zGaEOsPFX3i8PeKizOPB3sIb2CZz5Qe0iBDFLy28JJtDplssiaakFDKYfMHxwswjd
vBlpGFxCnjJrk0N/fDatBe8bxS3A1x9VnxBGWabUPbV5Xjjcb/NX24xe61yiqLJNNm0oYqZjZqht
CDpLFC9WzIasAr/ku9nD+cVeOaQZvvLwolPrKIdTKdKd2DYIkP7eYWc0h8stTkm/9paXqLGQZRyp
UNQN6YMBNmvcFCJrDnWWj9KXN9K/oRCJBt4Lb38jGkUxzrlMSOvmZ6YgqUy1ogdWFXGnssLIEFTP
6fjYG7GDe57AV/Y+paIj0iqFdMph+SXOSlsChfzNUX/sHH3C8ewSpJZYD9bEjQNoE/AvVDvp4uSe
2m4g/8hLgYmGJUOgiuPVyT/BOyLWg2GKzqKi8fsMzIves+qDZA1lmMSs0v+rG6JT2Bgj06ee7hsy
hbpjA/LbfUb/HH8DqURmWhmyw3cTQYQFYbp1SvTNL7yFVAP7J5aad1Rw3T86ta+SmaOylic85Nms
w6Sfrcqoik1G0B42yeYj5qE8rVZLbre+Gplak4tPkCv7n00Ky6PA5hgqkLijbXvEtXk3TxYHg2xq
k9hYaFaeSa19hFFlB3/2PTq1sQ6f0VEgV5NKHDZw+lC1xPqloqZ8lZtYHr+BAj0tVOD3wqPyHvq/
uN/eVeYIKb5w23bIqMOmhXNVUw/KIWMDx22DQQe88/uUFL7ZtwPkOmShSnpnLZyhlwoWroeqaEBC
gOD693yoetiSa2eRTtYhC9AmPXgnHJIyNdFlqoTjD2wWqUHGNrKSLEjBXivD00ZxIjbjNLAQh2EG
XhjEyQAGhsx2xO3Y6oU030cQzCgTK70T7jpG3efV4xKOpfqHHPx3uWu+0v5hyGE/DP6q0MQ4tcW3
b1++FGphcDAyB6UOxCtdUHBQk9NfFwbdLEAv0oNQcPW97BhIob+y4H9dZGLWDk3nN+3NnN7Z3Tc0
4ghtsCcn/yczfcxj60XuG0PtvmPwOq+l+XAeQoZAJxNdQjXqa+e8IaOFn+WT9nYbk2pVmZCMCkFV
PWfhMljlxhR73nCOPwdoiHo7rcWZeyvBNKIPz+FYWKVcWMLPWSePaCQRvRPbjL4JIxTksOY5OZqp
tzaJXU+9BbSDXOl/hYkg1jfycsIrA1HzZEqLZCWOoBV8almrl675aotmXgRzRLzOMMbMDoC9rmmd
yPeqEmqDX+jYAkShh7uKO+gOybVqkewkffyLosEwpyTC745nUT5g+2X5WJvmTKpLIMJf7dFYwsNt
dIgeFgP9DR/cRChVEHu/nYt2SdNSp831TIOotWb4KJM36BzXxKEEogUVTm0mGZ1QTQ76tQW5A94r
fSivokxirOxWj60U+ah/OPfR+tFRo+0Nb/BlNLilr7SATScmg4NUeGrbfSlchHvloc3A+sTPaGmz
+ptE/tedAcuFxR2S1Z1sxXxerljPKdz0qz0GxCY0R2PwMo7pa2UaiOMZci+kU7fpvOP8JXJVONl5
RvVs9vABlW46atBZZ/f7/wyPoWiP2XHKCRKrcwJxju25GPQDDsdY7sLDuIoGuLi8Jtx0zN/pbF3+
a9Usb4AhppdbkoKT10BsSFNk8m+MuJETU0GIKS4Y93m49ameUui8CmzUOtNTnp+f304BBOaP+fPE
mfBWUHuKZNTtTvCRIkIXaoABVhhaRR/LvzVd4yUsggwhWFiwfksLG7Mv44/8XwAZnN7Xv3v+cUvc
SFxczXOMypprWyGtgGnL4UIeF+RNabe7H/PLemcIDE8dMMH+LK8K9Nw3ajAWNzTYZkGOKFA/QyOS
uaH/9OBTT+g4LnFpjUALhwO5TxkcNFFII6Eh9sJpSdRaVcDV9CQB1L5JUxNarVL2H8iHwEKHTDH3
sLg08kgyQ6tlQufsiWbIR2cJ+2HNMtJFeXQXKgwj8DgJM5nzUui5QhgaM3BJvt2rJuoIlfYyhAuP
RysMf9IueTGBxUN5C+XjxKHiPX9kBGX6NJD27tuQHAURab5L1cWQNIiLNGCzVTHMOZ4g9SGRWkUE
pOdCkuCWYtOfFXRDyfuG16Qg0RABe5g8/UlpCJiPG8rpFW7BFOM6n69zt5zcwxWLGesQf7LMCi6w
f4+yqZrf7DfBfRXmOeZCaGXBZFG1tR7sZaEjKqHt3EFTMdmY8CpI6LLr87O9ByOV3WBIQnEhlcbu
jqmFUPhTWMFWlUmHMlFjSyyLQKQcHIwDi+GqWOZ2h9XR/peV0MkSd+h2u2QI2+DFVz/c31tVYkMc
YnqWn31/K3Q1nFODv73/ujQHmtpYB7CWiQRSFkIDCNsrmCDd1S1pduVJCqmH+5AbaKwKdb1MpPU0
ESw2ziInDNjIA93jx3QG7H5D+vUPmPUViC3MqRrx1G1w9/u4CLQ6cJait7P80+fdgw0e90+IQ7qE
+r/hV7ZIWzF9DTCLVHXQpTqwrbRKSB5h6hM9+5J8qA5ze00KFMmU+VEvWDAoEApKD81zI52PkEVW
Wx2cwpmJhqVD7f5sS/Fk3uDOvxM8P62efjdQNrfTxV4t6p14/9522kIDKKkhpWx72lftqtnfj5wt
6Hxr9tjzoFqFnDK7ON9AGZK8RjUR7spxF/sfs6VrffMZ4wHrRcQXuSUel/F1n0Lq8oUJ2/2bDfqO
cOm8q/0EBAxaOPZXoscatrFu/MsUdtAYkPbwtGSX50aeO62fIYoU49rJu8dwATdnKRRj2bcavQbl
j7Kp1WPCEGEq9e8Hi9hozGPziLdude51yhMvyAPsnrX0wKRi97RkYMaN+26qeqgb6iOU+7NaEhDr
lmGCIenyX1vZEFFUUAAs8Hi8na6lieSH+0p34a4mL42HnZt0/RRMicynq1nHH4jgYKaXPocj93X5
ZeQZTP4dynUGxT++i+1RoO8CnKuPlxN0GnO0zE0YCQduCgSMXYz9a5BfQhH4Ux/1tlKKH5eEZ8Xd
h53tcZInspGlrs/ysRilFVIoTn2qGlWxfhFCrkwIVafyfEOEaQE0kzrDsqNmrtxaIXgzCOp66yOz
Dtcdhk6tpJ4ja2cBasBx/yykDp6WPzTnneaa4AK21pNnDHkv/u3yCpJNRLufdilombw+XX1heB9e
AK2RrfebGrY8Qgc9y3paBuvt1fcxi2Ep5RdqGB0aMEOk7s8ReMwQzcSgvNlhvQzODpUOGU75yn2Z
SgYiiF3b8a4U7Sn0LWPu8An6higeQIuMuI3+iLnxX8lw6Y1HsTimDWCrQ4aqg6wLYWXdczn7GF4n
M72L8ljLStxyi1NPhB2NIrvPWd2rZZaXwWscHHBseiFVjiaoT7IX2UgnlgJW4z1VP/Wq9IIbmvMF
MvpLMVrhCrzwDyrdNVehKYMRVS4BHlmsCZvCAaZnRNgOi+2cvNlwM2sDxWaQ+M1QK++G8voDTPpw
W/cO6tkKfofAasFYNWX+Mhc4al71KS3SUq0ucMEUWiDbTtaVu66i+7sTQVuSSFtcJwJT/hYdsRTa
8dI7JIEgTSxgTVjjQszzFmbCohtrrNENvFKJFXAMdv30fZdLvr95O0Kem3lHStkV2bLMOSPpFlvh
C+1s0xs4Fvb4YdOT3T+eTV38oa78425A0dyi2MXe1fNBG/ZZbsEzGBb7EiJ0pO8K2g8qbRydcQIo
Em6Kc3jypRPkpSBYLj9cKMsOv4lL775swGgMS7N3zsEOwLPWn5a7yF4iJfVKuqLbaSUKxw57m1fH
A7Za4ZfEatNEoFnjB3wDShITdyG8jTG33CfHjP92aTep/u3fZ0xeDeNb0lKp6gj5IyJ2G0xwDx9M
oVsgCkeK67SThNIYPM3HYvBF34XUNytNKlVuPZglR6l/whT5QfDaqfIUFk0W2n8u+dKbSv5uar3Y
y/pKlWO6/8wLkmRGRw+l3cjFMFP4y5HbgGvYgeauam/AoIbFu61v7uT4BlWBJOOtmsxX1NJLgGhQ
Tk0e6/s8l2PX/r9tFDgLapMTTYClATw15+MqQTB4oJQK9w828rL7Df9eYUjYLAgNneioylmds3J2
fzPuL/maYx5uphsoMjlhi8xD06VlVv1kYHLh0Gvh0U/s1G06Djorz382LwLmhMbYCDU3YVUONono
2zwxYqAWoiSe3BCtn0Xx8UDyeqWc5zchr9rqPGR6k/r+NI/E7YmPvWzK/Hq7DlYqqnCQJEjWRcT7
vSFr3rn4OgHe+8OzVAUzYKhMuXxa7qNzuwgDu7NQsQWqnR57HL4kIXQnb0ShzMC2xHZBdP3QKyfK
qABt8FuFKoMKSwu4odynVqjOP7x2E4FxC1yV1/vV7WisLoMX5slDsxtWuZZddWC13+kJU+mLCBn4
Nhaz39zfPVERmkHrpIB2xTRAZYnLknD8gW9prN9/r1uu1yYYp6Fkw9+tp3wxETIYRhfFSab6Sc+a
ZHRyrqxSZr685WZQ2rq88lwEJpk1hwl4eXft5E8NlpopKOPTMjsgDnxSM/ohsWmu2qABKGusWcLD
h7ETQjXWDrr9UmhInzhhayLzqgt6yJKp1CUVftAO9ZTB8+Ma7gOCRpPJHR04xgWTrKACcIPn7mWe
9CyXr1rnmzOdvZHhR8hGHXwUg5NXqKbGFLdpNUbd+TntrJQwM98A6uQ4WNF3GDz65/iHyKeJdwvS
xsC0V1ymwc9Gkal/xcMigOFDq0sEvpoMiS91nR/P2pkq3R0tOC7QgyC+f9EahECS5H8WUt3O9naE
T+82O3SJsZbaaoeNl480Ql2RR0G6RvwZzduirc6CV20ZdR3AFSUHsQ/oXza6PNnh47LzqkjTVp/W
CnR5ETNoskj7u8YN8u1uqUwGq8YQBLkHgXIsJHvJsO2ObkQhle2TGQ8/2CW8UvnyQ+yJsAkRd4CF
0hhpxBOH3g0LmTQHqNgSion8/9i9L4ou9p/WhI00wPy2s2pjQ7JqeId3Z+RXzKtQoxVEeOg2nzDR
4/hzZwfaUexpsU3Zm74xg8CjBebqC+lSkQd3VTsSSnJpZL/8HHVQG5g9rRhnIGnuns6Fel0kjV14
vmT3pkKbXykNQlmB4bOjt1K+pVIsTKPxP9am3iIKzUN4cgnmnz7G/jkj9QH8A53pgyfoWvu6HUq7
TUfmtvpduhERcWRYNmufLFC+paqZ+qbHXg52pbZg5TE3UGn+psGhhq+y8XRcdN+h5yzPPZUf5zo3
pNSkkVKGH54/AMaYnvSZL/aXLNMGduPRqGVkw5/U3UwCBDgC8VqkzhCz96ePRelHc0cSkJSHyExW
7Xk+PodTg+Dpr8LjzutHoE6Y66HtpkIo0daS85ZpNikIg1tBemiOrZ6LWEcxlrZSHp3zELoE3vKp
c5Hw9onXY78ZChPrvIh0LZW3zja50EE+QLyZfPeAdNkaJ4Wctc57fkvZKMpPVndePV0Ko4s767lh
OO8E69e11XnzckPc2sDVwl0iFWE3WUMJw8YC+2CRFrhgCxTNUozoipqOQXFJPZ7jhkc9kcuWhPWz
HZQrMxqDP9dtLX3CHujhzeYBJ7q5QYVJU2IJuv+Nc0JjZpsMVYiMVjr41709ZkBkd45N4D7jz0HJ
zWrO5xVFjzOPKVB05K10XyEq7QFhX5oaSrcUQ+eVUaDNodt6Erx55jvN9b4ffoQyNZ0pXL6T+85y
hAiz2IFEp1+JEnQeA1wDRC6I5fXvv9wMTO4VYwavNyhknRy3ZADejyLH/yEVGPxtJzP5dfGyHDGa
/mZ8FO3FPMwQ6pXif7B+abbZTJn3pvdnC/wLYvCTyvqAOlKbFL0VEFCIfkuqASVZhC6awwy3x77Y
YTMxQX2df6uBSVysCP7ICWtB1/eWY9mbwktXcD/5dKZi3m7UUOfJvn5LdKF82auXtCHd68i84gGz
pF6ZWaO0VTb5OvYXjft94u30kxCRB1HEe/YIujfFegcI0mVY6qDpRk5BJtX4O9mKTdGP63WJsEnU
kt1DkPVBzUbbE0eqS7SzGoybO+VTfcB5xdEPubLFuKvZKC0JfOzrmbAMs2quxaJ43ibM6gyBQPyc
xGqigGwCt1HoPoQoqnuZzx1aDpYAKKcpRHDERb8oQa4EWPuTYMdVb2R3LVaT4zf8twHb1HHqtIA0
T4byfowb2HWNbrkjiL7TJloBr53GL3U0LiUvNuQD8vfms5qqJj5AMH7cjfboRG20J1HVJBdp8/Pw
3AUaGTvlkjklQZ6pIQINTNFGrCRfOI5nGV9eyJ2rFv55b8HrRxV19tYVxS1JdvJillDQG20Png+o
/e+Riz619njvYshRL+8veQxokZ4ms2Z2rWkRC8xiGgRE3frS8HmZa6sUAGPxWENqEddNdxRmrU09
23yzYKcGn0+BrST5eFGJdNjUOmZyee20v4axMw09hPF0x8DAXqN6kTrHHVUXV429Um/vMGUEFT5C
pM0gb5YR5fmA2b6GGUaaLQVY0Flz177yeo5MD8Keo7RfhpSFtaqYZVx7F/NxzzplGRxkwceyRdEB
FLbfI9BsTm+PJYUqU8LaxXzxfrfzjXMJ1QyHi1GMJT8QoVV7AoZzJs4wO4jKEOICKIq14E6QsXAg
ZqVzIrF4tFqhBNkCKdz2R/9vxfU0t0KPvVLo1R55G/YRYjbVpJK1725lM7Pe3ZesFCg0J3V4V6uB
r4yLgWqIogWYVwRXVD3yNUq4Im5W06NfyQla7mmcDYPfTpjkYgSabt62UbnUXuMNZ2L+a3dDrM7E
M7CK0Rm58nEKCkR3hNueAyhIhzg8ZefrgZfwrjYTvxQLU9py4UpGJ8GaCQzA+NV8C+n1OJHvNYc4
zAmORYILHXqNOPnSlLYxq3hoBdQ1N4zsA+emAGZtkiScZpTq1IEX3qcuPVx7ZFyoKYxhzJumL6Jd
dDUrRNYBNKD2YmJ+lUnclnPHojk4SUVg3GMGnuTn5C0D9jEaKMoTZGs6OBfVNdoXNeReiKH2L8gh
6sQxa6LPlZ9Z6cX+WcaQR9UEjK2XS9rIYDyMwAobfwzIu4n/j/qFfhDFoKvvpSDWFnPiTMLXI9kK
pGpsMu3z4Ihs4ltNyBuAqo269LLHDLQl9cwCZW57I9ux2DuL+zv5y3NZBDu06PRvSDzxKjd8925A
hWiTF1KNlEr2pT9GrI1P8Y3ODNY/WyMr8Jyed8pqlU1OjUssAEbuz/g9xZre6sydC9xivhyDYkP0
3ww6ZCqdTzQb6Uj4JUqY/+6ZKbYeF+ffuKxhI6qZtZqa/LIIJGOoKN/qOgRPK+LjZkTdqvfyh5Zg
ovBekfgbPq9G/GHGG4u9Us5LbaIIIpMF+nj3dHPdXrByMZZgp9UOlQvGubgYbR+k/79rlD+1x4VJ
cvL3HgenI8+sN/G4smRAFVrQuhTS7aoLk5NS12NqJS1u+Yt0gbnEQlg8Iw6y39wFzL0oPNTk0DrL
E2u5Nb6FEhpfb/NSAC3S8ahedjq7sZ7JyhluIciUxpFiUP+kU4bFeFyWh+CeAPfOwfN/p/+zdKDR
i4NkkHoHQlyxUfqBzujblP7qusS2IC5OZUyJmrDSdkKcsktRap9drHT+0QDFoA95APN8Z1PjbauV
N4kQY+091nZWO0JFLY/cII8fZRqiAUmLkC+zEZMT0MiWYPKX6cyOsXlCY0aUKeh0j4TCpshNfyHB
mvwr3QN9ajn7m4xjFHdVWexPklWLFfAnQTMLkVzjb7YhvMe5aYK1iChYzcMr9Gz70lQvXsfJt1Kf
QqcFYUtqwbAEUfA2aIoi0TV8+wXS0/MkZdLf/143d1J8x5dSY7MS42n32ZWNQNdJUZiHZHRF6USV
xGbR81RPRAwQf+Ag8wIaHtVS8H/djjtGwStw6CpJTwxFn8a7zoYJCwFAt6ZCdzr4LKNPN7oyP6zd
mv1ceU7ITzYZXLpwCGPZZ4V9A0zM8aDcQCn/nk/BHXGq12Rn8g6CsilRVKPgJ6W78FbgWCsZKx2j
PTe5/2Rt3sVbJx8Bn+CtmJHO4hXulPj2v8K5xWmdYtIWAfWLEPDR78sSIOHh+55INYwODmhioq0d
tWtSmSOnOt8IX6sFqpkxnfTX6HAMeHAQzkg3NJhFc6nnxqxJV3rDC5Crpx81YrX8ofwIoVyrhhlW
aiJ0sREHCOFbfNChnTQAWsig+7B+K5gzufR6ikM+gA1ShObvmoNa7DyURRWzXhtbHVBNgTlqiQsO
MydgJ3DrZN3ITHcOP/gh8UpLtZ/mVravUIF8Lq8sAVugC7FghcA/+CtNXtaIvaUQU9SJErFOz6X2
J9+BcAt39cMlQQWP72VQ2d/bF02FB88eGHL6kdHC+ZZlxKbp9CKkwBANaC8A8mbyHyBNXJGMkW8j
/18pI3Xh3WL0rr2irwowGNI6t6vcDB3Yf02dnoPTzECOyCjoA1KbjxSl1x33PJaVrn7zlI7zv3gw
Vq/kfzvneNK1/X6NoNljZjGI3c+LDB6PYxjrYha3pPmj4Sdeqax5bGxpt0d2qY7cWhTa1gAjDyvW
cbWiKPVsQ4ED3x0nC6X+nO79eR5+jCr4lvBhPW4QPdSyepK1yvsnnSGewCNTTTMWyOT4cJOgia6G
Md0G2cOOA4Hfa9PB8zlWXnCiHCRiT4JQVDfyzAsTozLcbQ+XCGmzGOKUG7e6ANmH0cYGMGjv2iag
ssCosicpwL6GMEFYxC4TAQN5Pf95mRd8P0jsTOWYKwlqidV2S5ULckBrEHBkxuwIPIWvncYUP+gt
oHvo2eMbkRonhQ0YJnIfrUTuLISepEWFcg+KeYuWRbXJ7J50m5Qw5LWMDrWNkOzqTZCXIuRugGss
nmYSe4u2zTAu9O/zBBLOmLdnBtGTwdmfEDy+/68ArYR+WLUgOthUX+I4iiVwqop1VQu7t2fAk7Rh
eKxZpd1wG8JJ9yws52u7tv1GTPuCHvCn5rNlONfXEpjx9HbPscYEv33HS9h6cDkxcZ2BI1oDF7bk
b5eEOt81bhZOH8TC2b7/wLMz67YPc//Ay5hGL7cuBeNr1QAGWrFbknkhOLCEgTUlVU9dBB4NwiMk
xImR8d8a4G2W5ECGzN2LyVz6ePjqZbni8Vy9AzznYZYttRq7iImefpUXz6EayiVGJQLLimRdQGs8
pZMT6yLZXMdCRvNeX/5HsjTHNRQ+rodhCBNnMVzmxxvNAAgDRM+t9DOU1U7XmI5qpyQh0vCNq3ks
5Fs2bMJSgOd4MjWRzxMLk0c/2g9ZYKG0aYHPkT1VG2Ly7ui4beBPuL0kHPumOxiGTeHkhxs7NFMt
Aa+RnJFza+bkI7jtrrbjnrp0bA7h3nVHo6Y9FoF0WoqH9xIRYqz65T4UVSuqZ0WdvL672GrBzPSb
ZJIzEH/iEzysMZVwAcaLQYl/P4CPeOCmnAsPqJMuACQseQrvZMi3skGqIBD+7LTU7e+KUJa/ThY3
7A2Y2PgtHDzpzmh5ewj+iWVgzE5lC8re3NTQeAT/xLCbwjKNsirRqbtJGZg6cmiX7P2EZOP4JmJ8
MAhORdIdBN0Fn946hoWbxdLdPxl/EZqx7ftdyjZvICWueXg9nAvZ9DL3whfOfJdMWs3IoYu2SHno
mlx7mxMtAzgnoTkQ65GRIMWpc7YzqHtBBEB18Kl+dM6y52/ISqwfzOqWOkCAYuTbmR3bNCgC8YjI
Jb4Q8vsdZ2t+1VKd4XPV6vggt8q3bIpRwn9iQ3usfAAHXbacWUl4N+OeUtKUeTOPaJLxCS2vR7nq
waHpmnMNJOl8Hq50jT4iqz1P/u5IMJVQuycqJfcbwBY6CVJHeyxUgg6SDtPlYrx8aKLAkL90PWy8
Sd96yfncWcDpV1iQ7yYpI+NdSpOBVdVHglLREXp7BRmIRfUJWkf5+6ywqgU/I5I8NoN1n+07CdIB
38P1TKTjEJWu80PA3Opt2OCV8J2Kji+787qUEgsCMw4gpfnQhP7A3qnTWHZa5JfknsMzr1NHFaRx
4qrRkgtC87jJ0knY3+ELIRwy944grYBQ87dNlL0S2sGYruyn80j1VTHCFymoVDt2sARXwO5IzJAG
x8X8TfOnYTRGJJ3Cv2PnPD87NQxq131EvLJg94zK8UBAogeO111ysg39Yeg485Gl5goePhoD79kz
csS0XUkZGnIorrN9nOseFSQy1EOtkz8cFrA7HySBiErk4BtHi7QG+G9BBDeFnXCLJuQZ6dScqEYi
IhKey4tljYNQm+ptSsUXh9AIzgxwmmksFHfHK5YxH0PIC0dZTwD7SdUTMhEypWGlL9UDFfFXB+Vz
7xXj9TaEPbZXgqrzxo71OdQeURD3LDPs7WPwPCNcoLTAXAAA+0PDhD5ZWwglMax5dpc40kHu0uc8
RdxkWTATUffFVhmQMvU6+f7WkU8xQNTz8oWht/3/ECdz3DnbwR4Iwbqracl81ibHV57iNHGoXWQF
yigldGh9DWrzEbRMN4TuQrxXobZ7kFXE43bwVkpizhgt3jEGCq10V08Qm8Wgn8ag31CS947SnF0W
ckfuPUnASdcMxFRkVrArcszGUEbh4G7dVyUXPu2lojooem4Qgk/d5zUelw4UZYg++qkyzMDYRYJS
MuUbrp5Kl1OZHSafvyY3RL64vmYf0GVj5z726k3rjpJFaFvTwORlET1Nx5EYN3eL45I4YU79/3np
i8OJvlNSkdyK6nP9NljSkshj0YIkEKkJyczAad90H2UatGgJZoEBch/OYkXoXwFDGsbJk+PVTyRt
bcpZZY0om3itHTPodQar1qRS9R9DN7FhfIo8ZfdfmRHg/vEmlp3IcGPuL8COEPmnP9b424tpMCw9
SRe/X9+ff/LjZsq5u7c1CjDc/zvr7Rx0hjBYvav4EPpw0G3MQaZyqy9Q95S3QfLEvVv9YVbPudZk
7/RqlOcuAyr+zBwLzDDGvqYPdpxNZGtnZP6i8CqoXQd5CO1j4/DXLuKRVDbT/OWAKtKeU+dPqi+r
AB61h66TOd99in9A2o2DEJ6q6rAQDHRDeWoGBAvgdACw46C6QDvDreBEcdm/USv0AwDiYdNxfMZ2
tJt/PsmXRuhSqhqWesMZ/I3KUNu0Hto6PF0Grtl8GDBk8b3W3cq3ao/P3aVi+bNfPJTu6ayUGFvW
2VkA5/TrU723LnhMINjG4wsU6s5jU6kHxBsCE2yThvGisU+taYBrKH3AUjM9SFwUhmHpovHmAlT0
mv8CoT5tsrdC51UDnnQJ+M4iIXwcuDMNCJ66FgPyAl2SXl3XslcOHxZWChcQEp2evGEkJ+5s5Zug
VOoE9+Bim+9Ac1BtMiTk9LjLJyVJh1bC7arSgzcnDYba4nbZcuQXVB06ihAW4iBJRlmp+zujORKa
VqDodKNuhEeXyBdjCncKDySNHz5rDU2veWo5aLZ0LrE8wbo4hnigvbzsM6JUaCVT5qlX3INE9ArI
OtEKu3/+viU6/uGJHH0hVWSCA8BuFfrExH2SaPg9BBpu+CRTdEJDEcTwAMfNi44bydzIw94KOi1O
E6RpcWcdo6YF2kU3I8vLdZ9j628TdzlK5tzeX07Qz/xIQdUHkqvp8DfkINbq3td7/ACvcIC/CoLK
/ZlQyNI54S1G0ZiXgzRa/5f6iRFtqKJOWnNf91Es4lNw9Tf6ADT8/a4GBvNJZKg59Vq0LpQhhKiY
ISqfvyzmWH8SnwEvf0MSEBxutkAbCsBGXGtO7wcvT70iszXkMbZZSyJaQoZtHGlThg9i1ls/5qmi
/gtv1Z/pINn1H+QoWElnq0qv5eUX11FRZVAo4IhqEmZaWv7OtRta/CLAt7bRBxgAa/R+87PV9+C8
rp+rEmcwOXRjI8trdIF89GTFuf8cEHQGu/Bf6Ioa+rcFbp9YmxsOUpIItL2pGZfppVQ1in4e9HcU
ej5e67KEmjfRTssIqUzNP4p/+TVCNu6F8Al3t6XZy94UJ46K3Kz3P58SSZkdqt7IO9xHf4zCVYjW
0HvFRlKwGc6JTYh7ZHg8EucOwEoCmchH2/Tg6QYaK1DAm1WyhqE5IEC347Wls1L3LswKL8QFPUe5
XanWJpkxVG5csoOAZkrs3/7xy+DY+qeb0PWhCZuMmwNFcspMHqUyL+M41w9daISpbGjS/0Ivv8g0
3xXUfILsHE91DVj27ooD2pSytwxakchLsDmr02EA0rZD0cvGV507PKIWHN+ln+XEKSDixD8+Ia3y
8cp52XytBnHDYm9izTBlHYR9wVuGgGoRpKSqk5YMgvm7oBacRc+DTbkHJ0o/BuHPHENP/aLzau42
/Xl8BbCyUdAz9uHrrM/vN1/BqhRp5EhrIFA3dNOW6iUrq17JLl95xIeLVM6WmXTAUdjOa/DZhlcu
yGNMfJBpZB7DxzWTPcVjqRPj2FTlVzqyQdiZu7hedf/Un9Msx8yevvLG8kFMPq1S2dnO1W0cVVmr
W+HShlAA9KKbwncCSTEmGgJebS5a3Nv+dk3HC0EDGRcRxzV4fVrF7AzHex7J1tn7cfexx3GosbXG
grXQ2XoEPCTgI+XEHCkLX38VeYIQj//Xd00n3mHzLYgh2N7/wkFBPCSu16kJw2rgcrNbmYWQd0OT
cCHDKLMj5oJP8r4BsobkSwnI3dm/3z+dJzxhNJe1kUBSb9J8A39zsbvkLzlz4HDZ02uWKWFLhNZt
7n4DJjB6vgUwfpjd30sVju5+ewbQ63zPWo/R+qKQQ8Y1x0eDYWNcllJSoxBSvRWfY7lHJ6RRCEtt
lxnv9YFLK6abkzEI+bi8MZCc8P/SjNrE8jc+hSUiswiwPY4WZNp/y7v7BYhZmkLQB1VO1DH2Cx80
JU+t1KEPx+CLhmdwSoIZgeEpnGIpCaR3TvKIFote6NjV31T3ax3EvwMjriBHBsi4508UUjYDsH4e
pkwEnRaVQ6N9JXVXAfIlqUTSH1qDsPZB/+nQxkyjYH2IBKiIuPUbb1JDEmDnfk8E0pXQhU8OEGAC
Y/Ip8dxJD7V2q/f3IpXDRaBM9ZUpLNY6mYlwKAR0nicROLk+1PJFrN/GtBXE3h8L0zYyKOltQJeM
89l8KENQawdPrG7XtpO9qXxuNHTDv5FNlwbiWu4lz98AEQ3N7GykhCTyuzieBPiOZLs2PYsutrjB
H44d562/tyqlPWSknKHpiwSRdCDW46R2Gvn+dK+73jhbPYNPfeKaUCuRz1eL2L7FawgvwD8DeWcT
afAoCfZ6I9RsCYdmiDXicM5XFUPDOjW5Ff5muZVBoraCYPrNir26K3htu6yy+Yhqd6c8YOFaV2sw
+nf6adyyBEDjgZGIuUrkZTs1eYNcQteWD9Q1qDGdt5/l85qlBupmzj2rCdX6JSK3oiMbAzYd0AWQ
Kv2GRhzx+4JOJfI7HVURlouEXZd9qCs5Hm6GDIWhB/3qA/kPYEdrVZiEwwRAu33FCqsAu4URqGQF
DI46z0psqFszz8WgXl1h9SNTzzXBKs7HAz9DWmwtUOWpn/JMviAQxFfMPlYwJP3AXewCZvcJbB4u
FFwQ1aqIGaC4ux2J47usShm6ZmPo4DE+x8hpGTNTqZkRMsqH6r0N8XLALHOiJtbY3EFWaHCMbSsL
nq4OjxqZX1MoQ+LSXnKgJBUHFPXZsAUClJn+DqnL7UbV4odZmz5NJ8ajsNw7dZeIskqwG0USymlw
i2iWAoWGNnIdCCvYcOYmxyMnUJii0pS6hljJ/qV3Na826rQrTBCV6gnAkVnKT+XO+S7B9NKtPJbn
22KRUocE1DkOEa0Da2mvGihKRUxKxZgZBnnJvlOK/h0M9o+FlJrCuBWLCv0+veSpo4GUt5pVh2LM
Xt0j8iX1mp2Hg3Cz8d5qlvSw9YjwLKTIyja3TOZ6DdiwkvJxjkJeKgZ37MEGl22x7qvGVKjKKhlM
vCBOQxJ3CC9l9AaQVIo3peW+FvgdL/ERHM8pjT2e6UPi283veA9NCp32mSwaW5CXRU82NsgYjAMB
FdQ/MKAPiGLh155DRz5ktDComvULdIgcueFqRdYJgjj/5u/ey4kTvqr0uD6Ye59J6EyL3XSC/X1w
XtIwg3WP5o736ZEChZVhvAwPLxtgcUhZFLvuxDkXsVw7UsRSsY6CQdN7qgdslgW08gwBfQkGyOoP
CkGP/tY1gvbO7MbGiWkhZxVEfT81xWyLyQQwRvQRkX6fn8w9bBvGO5rFpR7FkbiYYfhrMKIJL4UJ
tzo2nBk1jRnxErOG9pE5Dne0IYCgmgJ6RjJe9oCvMACjsmXHOHRW39quQSGHwezrdTVeCpEASD3i
GmK20K8H8emqbf6KLytB6Rv6P+dZnHz6kBblibQ5M+Mdwh+nT2RfT9jIvH8hiFIPwe95nEu+L5kn
9f6H8ReMjjRaB94dvIqYVIISdiq7tu/ZDQoKDYV9fswSUf0ZTF1gVi50ezJE1QDE4gqDXhxR/gmC
CzIZ1YfcCeuUKJX6lv8f1pcocXEYm4atoXUj6JV9gPs0Y0VmuyJOvl/Orrf42dFuk8+dYpPdhJA/
ZWl2DNvfFD+CfLyUDkkbDUSa+Y5DV7tbw7TiGCy7x6JKLO6ryyQzhOvfUm2/b0T/QvtvatCyTaDV
qvGYbuzkeoISdn+DYJLmGY6qa0+Y/NbgfLf2iJAMuuyQNBj8vi/GL346NxvUhHxMAXP3s7dq2wsL
G+Sb8KO3Qfi9WR9fiP3EQzFQ00XOGHCoYk0jlbSMe+EJfbBtEYnLEDV+uP13n9Q4ccSWWlXKu4vb
gqkEGu53rLPfJNSszPXrU2sIRJ4MzqigkRTc9eull+2Z45QCuFYhiimfZ2eYe4elcFBezVGqOqL1
1vsgLFCc68MvE94m4QLxk+psyjrSblh5XkxAQ0jTC8JnLvldn1GUcRPu/+V0lwpbqTubuElOm9qw
sK7V071dw2/tZ1R5pxJAdpGqakvpBZ+FjKTueNI1yeSeD+Z3BVd88+OgSvgtYaK3H5Pkf4LuhhGd
47QYHMX5Hn1Jj9+4/VY07X9GnLFHMeSGV1BHZ0HnHBfuDx/BuBwTMr8ubTeLpjpqHjH180Fxf0PO
jtZpd6PpPDDsa8jhCZ7cSAqg6Zeo/5cmF+a317eKNlDjAYU0msEr4SkeLXI7IxIQlTOwjkHOTvzX
uhjhqhJsc977Y9bV8Q/VAgIQIlxbSMrOQa8bgBnIcWp50HLIJCwR8zeRxiejXlH46ZWPzNGdU1aG
ucM5CaN/+A34f/8W5VGC/URhRJygR0KO/WJrvKaZQFkGJdWwP1Xy6JMiNe88N3/xvn7QQWuHKj77
aSg5AGN6iI5+JdWTgwM6tW7EcwjaiVU5z1mzwXDR/k5t2tMwd75A+ya+uPudqQ5qZzVCpq7mjSzA
r5MYsz0GPbrw0Ou8Sqpn9ld4S8EzeER8Tt4Taf1ox76650A3jn5DhElwXu/xrijWuDJ6d1AwEsAe
/Ym1p5Lg/g3rrPjDB4MSvGN2OiuONGx4Lvl6DkafFt1FTX5uiNCvY8MEoWVGD5vFREQ6xxGAyVEX
jkmBAbaCoAnxKzoXyeRWSGj1Lf5VPdofbcFPlV4lATa14cRqsT9Xp3uhBLR/+SjNlydv4aRS1ob0
ADTJsWQtGsPZ1/qHInpDoQVA0W/Ou9uqC/h9/HMgzg6ewT7FaEm/MKcC2KKkpjog5MNkPiPB4oIC
q/5k5KGCFO9vzNJ8OVeYruJCHK5xXtm1Y6h0i6OQXE2+c/JiHuYYa9wkA6fu2Tj1aoqPcc/i6brE
82eP6GJF+0nwcLIQNFVf6wOdnfnKsEovxOFnLqLpb31QYInu7+ZhzT7Gg6jP0kqBXq52++wwLTBI
V318HafuFm3/VoQfDuM4u73rpNDwGW0gRxvFyL4/stPwgrXIvMJrIIkArOF9GuJE3JK4KTCdzw0e
8sQmQr1d2p4erobaEWLdj3otI3hlhCgwo8PHPjJ3gSPeW+n0YsYXqqsx/yNJkkoeJyI2Rh96OCEk
5KvW1BXxPDqpMw1Bs2fSfemFQtCAi+zb344OuQE92oreVHYqiGKF8XIsTA2zS6UblZpD9rzQNz0Z
miUQbJNqi1PniUFtowlwCIYzAPW6hS1Mg4f9ZglNvKaOIy+1cHVOARYLGtvCc/HD/GJp2c8pTMQv
CYagryalcg9SaEpWX+7ggt5oPTjjpODgp+yz+TwJO2d4jSKFJw/sxtemd6OBqksr6/HIYqe+27B4
wMHcQGXgFrffQUcCiO78nY796Ax80YH0wDDQsx0Og6/bJAeVNHrCCgUZbDVwqOB3kvg0dQzqAUhx
K07HCnRcdDS0OGdPJTdbpYj1mW/JX0u339vraSGIWsYG1PxXHw5FA/3t1PSCvqv1Yo13CCw43r72
ItNez0lr3KRPG0+lo/wqRnoPlWW4sWviC39YhIjEUYfSy3OwkNDCCE3tZucJK4uHg1yCGDr+ommm
ZtAbVExi8qu4Va9mNj7SXB5thNXKk8qSAxQF6RmNL8AD5qmw62Jk+jKG0rYI4tfxxuv9W3TpcTgr
pfSfHKEu3qLkM9UmDdUQlKYosvPtgW671A8D6JSmq/LXchYx/mzlp5M4JyD2HcJ7OVba5vcZYErS
RzTeHWR2nGRBUpumFC0X8dYlzeDATbb+rGfmqBuMqE8Xlbkvd+FMwLLNdSP2vMAcQ6SvlWIlXV3l
Ke5SQrUE/Z3iQnZ3j3IxvYjQd43au5nL7BI7eKQBvY+R23n3NDZRxHoSjGxVLMIkm3/F3wSgVGcL
E6DA5emsRjgPY+X73+BK2fFFhwgDn2aUb0GMGjyobWIzFoE8rlqDxOCDo2TKqVWXeCGuFG6mUKko
6Pb2ogTu+PhEs5GK/VjNjgGsVVORfh+JTiKuT6FFbIG8TjcGE7AD0CbQfJa3f+5R2RbNLrqJEgkM
w7SeQAdQvkKo9gpy0ls7tRXRvqThtffLu5UMLgUY9x0roadrhQcicYsUYWUlmlqz1ap/M3/GLJX0
aNU1yey+jYFR0WErbN1wUROaxx0jDn8SEsKYJkSEONa5YJl5azR0VUfsSk3ZKV5VHYyeMy2flcLQ
4pa83JDlX5W8RB35jSnHgiQY5zu2yzCcAJalKW3mTWGEqeKZEd/v7MVKcU5xXVM8hJL8JXRbou2a
nv6l4l1FpM4OP+tCPs5+jf4Dxbf3vn2OGimZ40CS+VuG+BYRqjsydIzlpibzhDzBUGrnd0XWIVjN
nTo9nJaavlLh3X7+kk9rYjFnPo1ev+ot/Dx9Pwr909JSnoV6eRYxoFlsuf10/b33INjztpKD3E0g
/71X8dOduK2vPsi/ge4LQ2a/BfCij6aHqG7uD7ty+JFh9F0tPDXtByv0XNaW3UGzIl8LL8mjIdAn
//2ADskT/B/jyFT0KHUVNbwtTfMU6IhzbBuvaxbJZMlUGY7Af/HxTJ3JVD4vWC07TH6QHzG6pcCb
MrJxfeQ//QmWzy9NnnkP/zwN4jKNR5ABK/io7ANG59djx/Tsa9m84kiVI9FSiK2kE6rGctOdcLG6
TN21SIGRyeILQWOeSYn03VHLr1uKvGmwNlFHLx4gffyCeRcApAMI1jH8ADfPwalDsbt1dqWG/WCj
QvnmOjsipxlalCK5T10+tviXl0Sl8GvE0/crqxl9/H3dOAULagKZ4u/nDDR+J8RFnZRMZwQRyMl3
qzAXyipxfb2aZRQHTZU+YW/9GDWaRZCkT2DKOsxXOcb1X7hv8w2tZHT1BGo1YBJBrd8TS60FDPWv
i8mRO4h+nnA4ubLtEmd4Cy4NW2Fphb82gTqY/GM5sO0filPIBNTIOLRp0HDOZVDOVIE6HoxhFZFO
YBn7KOLd6WkKAJtJCgn5yYSUJt5o7IaDojNY7tCDnQiZURfe3jgBImwdICKXpjPKKkOvjVRwTG9p
gPaSFdsY8Ye2RiedZCr3UoQmgGWVkRqgWejz/VxYhYiMUQ7Q8q/pH2nY/BfUWPtK76J/jHtDpz/o
Sc8hlrFf+8FjNLIPB1IHVvigz+GbcD341sA9qbA1CI4pdZ+sBg4sk8Z2a+b1h1RJSl/Pg3azDk1E
mDPeYXysXQ9v38tueIyR5SBl52eDJw4y6hUxiRYjqLaUiObJgjnZLF+ZbQUD/513pp+zxLdq94my
3BkMw9PqW0/v0XMNyBIFW/BSghzUABa0Q6Jvb39WT3Mw6fPHBvGnPRTZQdp9hbljE6E9YYPWx6sC
4G56jBba/ozZsr7kOs4qYSFgTkVkPFJ34E1vDfSTxAfkYPRdrdNVnmdVZV+BZUNdsvFRpv/AAbv3
s4wuuEYYviAS0yCiaK9xNTI9IxrBq4lWNs5E70SNG4lW8/AzuCdPq5fd+GYpqQBCe0gPFbKYShBC
0gVRDeE9mXLFu5yiK7k49IA/Siq5MIMJTqEGdwWLpSshBWaG1V0Bw++DrF+QN5R7DR9CpFptPkxP
U9Xf0J68aIQLVL/l1Qqf6cDcyvkvMaI8n4XQMOr1Y9sWt72PiH42VKlwGcP8ZNvajgsUe5lsl7r7
y+G9FrSs5v6wmSNGXIcdIcDosysyYtyoLLUKXeyDpnhy+f3Ov8v5PA4MQGLKAFRcECChi9z2T2zC
v3fBc44GBGH4+kMhpetXNwxPJ93w4wEHxgi8NktqSxjsC5BXhVGqcnowfOiUJXUr9NZMigU5QOP+
64cwrwRA8WJfUyFCd584XrMDDqgpjHmgk3kuFqnXd5M3Dv8AyoSSLoztLFZEtuA/llppE+6LR0Bi
QrJlcDuZZjitlAo5gSl0u6inWqkmb8cAKEP05vXj+2qaHqITrpzeVdmyWC5NdX590JDzjnaSwHq1
3TmjJEQnpy90kF5OP7UTUqhjYPeoC7AYm2IoU00NeQIEzk8T7QUhNT3YTz3oLWdOl20XcWgz1o50
9wF7nWx4kzhndo0S9v8RKHGItGks6hnAHX7Gzl3fVF4i831th/OHv04lr3q1aP7Sh7tafE3W5Atr
UhJgCpsPtLZQtF1CKMO7m8G+/djeOuBoQ4UwXW+Hb7SDTsz3w747uWTnJm1+MhiidiL9Fqy0EMVv
e9EiN5XywoYXKHB+HPWaba20L9Ygl0rPX+ym3Aym/dvIHScAV2wkkLUM9rMV4ZLcsCOktdsEi5g/
oIPdqSOYcpQTzwVJA7PNmTQxWRnjjNRwMOm8JtZD0jsAMfMF2SgTK0r6uEsIGDxqm3jOxWmERoO0
lv9a9h4nwnPkuhYhH/Sdn4fI3X+sn74Hun1z23EOAUHZzeHhjQugGnAnIN/YE7MvpxkU0stunrMr
RPgMjDc3hxNhWqDL1qee+ADCucriiyvUzONKofCJ2OLMn1curO3Y/UJ1ck86ULJ6+7SDGSgwbBn+
BalxYwJS6K9lcnngrXcmgvPDCkbc40v0FzXywJZb2Jg28b9t9Nr03suERFZxfwHwbYqeWMjiKscq
XDInf8nILsAwz6rYmldqrzcJ4N2Qm29nlSL8emCq41dIwqUC/IGWL10qZeoPzpXTapamhsFjaFL7
+09pf+BwjHiG9Y+NocXsRz6uMEVSL+PglT59h0uTsBKvTzl/9OYmhBNG83L4nW1UKdt+y9k1pplP
tOSdyQbuMduhru222Y38MOFu8rNrFw4hHFRTqaeBAP7L5WkKAbbzLpqrTfpXUlXC0HROPWiXlWxR
o1ol3Eteh63dBn1YSyYdHgvm8DIKrEPVRk/RqPTK7rAu2LBfMbqY5MU5+zqz5wrLjNu1ixbh7vzD
4jhASW+29KEphLbq65vbSYIU1TyUm9AD3eyMrBI1s6k0PX9pUNkplMYfS9cVxYsAaaUQw/pOGHRQ
W5HxXnHQvMADp7E5tMth+/kzrCsi2/0oBEgFoTCMiE/W0DOmAkGsyvT0Kj2PHnexf8wm/jVpFqS+
6YZX/Fq01ByDuJf4HJY7le3rP4kxWsH8epTvIE2i3P8ZpvMsi2nI/8sB3B4IXu6Q82IJb7Oqnz3N
PGNMkUUSfvWiHi9kIgwJrBw8eCJ8K/yWHzGXngEeEG7l2iI96wlOPPb4Oi1CO5Zkv9/KQq4dxdtc
UZTaltd1Hk3IUll7dwMEzB2GqqRNrG8O9P+VZtF4/fCffYEgydEisPWpC/WS6Kf6wyqhOO/SyCKX
mhNhyMCdeg52QbZZ0ynSKgtRMFZvpQ+ICcbqDa+LIYZmlsr2pruQtlIw8XEPQZlhTzkVJk85exfM
q5wwMlh8L5M2OAqSDail1aPosDqwNy2rVfdFOs2zf4JFrKodycE9ONXhKzrPEqWBwdruuU0LZPPK
KAhxJ//10kHL0RGltsA+F6rD8hRq9QdkHDojFQCSRoTQHlq5Milq5iWtEZ+CzRZ5l4s+N02Va/2+
cWQL3+3L67oeC4Ekrnn1L9WmFv/d0EAX+J9APHHL6ewWxkyM06EsYEJcA8J2e8hR6CQlWlv2+YED
4PlUdAYUr4DheQ53Q1eNgmUVUqtG1J59bkMJRYdH71B1GqIBSykIu4QSZruNh6FTeP1KCYTLZQNR
HzJ7uFRdX78utZ8iZmBVBYyCUM0NptOWS59IJ6I+Qr88bt86IrrhXdwlyg6iemDe51TWclo4QVhd
S5hWGo4Bg49OTIeGfPujJ1bxWp5pHXUe0NxmuYw3RsGRb3IfPpaa+2n6Z3w3icCL9T13DbWwa/FQ
/ErEEU3GhZNLqqMO8bn3nD7wx49454GFbtXESett8DhjVoDfmtrmNbyUNl3CghlJ6ibcli6nWdmx
m8333SL1XIbn0xT3wPsdeHy3gFhgCAZIpKgiW0kiKMqMlVAfUr+zhIUq3Kcb9ffKNt2DoSmfrHwk
w0OQA9qrnNj3moiZSQs93ZsU0e96sL9VQOeXJfOK6olJpzYasOPWwQGvAHwfsz/S/36R8in/Bznc
I8xa9LBmRbc2mTW6W936WFgmOG/wmKcLCtSoNrVsCbwMEmizrx0ed9eX8lmDfBxzpPRJi5Qzk2xB
qZen7vak82YyD7NBZc71pb7IkqiG/IPeRXZQRpCu4oW+/PWA1kIvhNMtGHHDZLPCvPywNHh2u/g1
V4R6Al/4y8XV9o0U4UiL5bc23c1fvezdFFGJBViSHVjurlGWmd2O1dRKJHT0umfexcgFCW1oE0t9
rlNDmXFazoe2lbmd4yG5IN6BidMTbTsvJOHauVHLJpV2uW/dCqYoiSRR3a+Fx4gkMBqGaNa5jFmJ
exry48IPyZ58qzAXg/enQdFv98UgVXa9re/m2RKWvamB5Z9DjNE6TaWxYQRI3skrX7aIGv0qI5AW
Ma/FUm76+ewe5WNlRtJlZ+yP/Zu8HDN4FmL/pGVXDfuBM5hg32/oV7aHsYSJsGGrXVTtYoTFfcUq
DFFppo2njt9xx/bpNvK6wDV3useMqzg+a4+3zEO9cPRfxNSmtHNRbpVYjgFLT1byj8tVfr4mAK6I
AM4e+EZJVzWKehetxt07I9Wz6aGNqJcRXi36Wfh7YL4oDBv3rqFiaZ4vpK212lb7Ts8ZjvRA0nX7
laeLRkDm5cVBsKPWcBxwBtCuFrRvQWzrmKw/CRsAksDZjhN/+uNH5QG/5/WWoiCFWCvtXL1PRdRp
xX0CVcJZH7y0l5Qyll1wMmD5vPgGFJlolftlbLJH4bnwmJgs/BpgtrwIgUud5nGyq38WR0542NJM
gwFDtnxE6pkB7ESwMO3AddjEZmOh3E58uPe6oLabWsEcvB+nl4DksdHSC+wfXTlNXaMPsToIo2bW
zv1gOvz+mSiEbs9p6ldNn6VSAm2seIKWeoBTle5fVhzEueUy74bxWzM3r0A7urY2Tzcx2H12IDA0
9+/kypr91Aac3O6fCA7XKnyZYifNI9hG+UncENEVcldXOBYrt5cc5PmijTwnS86utwYcxiK5ceZl
LN1R+E6KA4Z7qtRvQD63/vZQnCNj2Yu/RwWGC+5WafMAbU6nyhMbRogPUICWK+jyzBQJklbtH5CZ
k095ZL9KZgEgDLMQome1QxA3UohMndWa6YoQka02ytKqj3fLkA3WUiI6BzESJY8IdU+d9Oz2TD6w
UkrslbyKPOkw620JCep54ugHW+mPmTL/Pi4PYSYvn/Jqy7ABzOKE4NABNmLjvZNJrSnUjg3BtHz4
U1ZOBKCG8j+1pzMN2/ct9nZaPRE0cfolDeJf1pozwNn9Bdb3S2+9h6ktvy5Kt6wZzxdufe9Poozu
B/12u6970U0w8XmqBkiCPUNiZPQXIVTo/tLpTOxB7LD0Z0kIaWN3Eeqwp2XSxauzyuZ3NQ74/Gju
2gf+3eSZ654sri2JNAxWMgaF98uxqnRcA0AsRZRPpo9CzLKM3wlJCwwEFj1iwKFzffFtReb/tWUI
VUHaF2EYpce8ZW7QPSsriDrYIgLuq2fgjgcsMHZ8vltp1yWt+bj7ZWecqD5hNwnwLiTeL6L/rZZt
28hlA7jpWjkSNt+ulaGjsmp2fJjxJvgjEYGm9uJA16LEjOFuRoq+8nQYgKsObWA+h95ZQau2qbrw
K/C011ayrvpl5FJPK51SmkP7w9M5+2E6Ypgjl7Lnmjr3QUVe8SISm++gNNZSSEfJsYOV3/O2LLs4
VzeeIu3hdsedjyRF4YV91iBqilsxnf7T1qJHlur+9hFwUgOMes+KODe3qgFZNmvnr1nc+VMi/j/r
Qc6lSqJgFREYHiFE3GcCFyWZ36D0ht4YFI2Nm2sQiCNDoWOe91wvuXxjdBo3H4Gt7+0q6ePWaWg4
ZHizkav96Ohp6u70D+HrSt6122V08rcPVyiZ//JcsgCHs2NzdrJA0LqEL43WdtNhHtjpko4B5md6
CBuhsyXG+kO4yRaW8wETq5A/v2gdzz0ELu/VsjNUH/G/37P4+E1cJh+f08ESlS25xs1Lrx/M5dLG
K2CExoAOTuR1mSzp5CWR7ekqUX6MNcvRx8aBMpDk5UYpRiPLb+tRpVDxJ++Qj8Y+QzqtLPKLp1xw
tpTFhg25cl2FXXEbbQ7CgwBAmx+N6aCO1Wl2i95ThsDSK/9ufyavmL2U7qfcnNZhZfKATeHk0VmJ
8APC3RbR4EWvfTIFXjoeGGDUDO4w4cjS0C6asEL1r/batov3ET/WIpsnYxLihSc+8js1kvyilhI+
OB1bFdyCnyL1SPxNA3PuMdyN20aZ+Ab/nrxj0l5xhHp4PwAD4lqqPy/yQlWHMz7DtO0FWSHrsUAw
d10NGquRikthaviNf0Wd5e9BYQeHZTCEitqnFYp1JGGmrTIGJ8hwruwgaKugrMZETvRRyAVDV5DT
eGx9yp4RQek5nttq0WmadxDWjT+zSx3/HUy65hE2bz6cLcHtQdmPed+uixYLL2fgcz5UooPhpPda
InpWv8cHXCITxZ0Qd3BLSp3ZDEz/l64JWglegnvTL0120A4P+xqdSX2wh8wo5HVBddP05xCuBzY+
CpA4TmcrypHcWqnAJ6rJSIdBnfbka9VXZ4L/N7FozMcEbX1ueDd+AUZLd0Pqpf6UrC03irsuvzLN
9CmfXExrmmziPu0aLtncBRTtfSR+r/IkpuSPHuBHpTSf3Iv9LipfelYyPIYPVmFE1LkhIcJNYOQH
QgM46VkFqlnXhW+QDvXpORzUJ1AzI9R80XvIDy9APWIWKz8QobJdhzhNk7DXPJXTdiDcmdB2lNug
b0po37NDpn9UECdBHv4pTBgRjCeU0P/7p1Pp7Q6HarEzbJhb6wVe1Kv4pYFw6klqY+OSJ7E3lqhR
RpPUngCHOQoxslXmQej0ihql+KUChTtBhWk7a4RuV2jk0bPkYkgk1WCrTdYtQDhmZyKYZxsQKEEh
7mbOj1yhoRr4RHRwaqBIM50uvp6BRlFeCn+9qHHHmXytcEoBUySi7672zP8Y28S0QGVkFk40kpjf
1TRFsHlwIwy28014PPRD1aUoED/z5MRXaVncCXErBVeOrgiKs5tH9mWsE6Bydtk79hm7NV/6TfKl
etF5uDabrvYJAVyX2S+mKBgDKglwF5HZUqQxx6RO5YeGHONWdhjbhtK0pmxRLv40NwMemcTXtdvw
tGhj2+ge9Wu3aFpIXf470JWVnkw8yTJbyLVBkPmC3h+BVusVuhdeifrV+DChASH0NQqY0el20PTs
G9pCc82fZF5bj3Lek7VGI1UCsFVjBTyTDvUdKmlCinsul7E2Gv0YBzyuv2JvGftT3Bft6YWQ+fhq
zjsu7U8ZXqxf/eVjMIdZ8FaqF1ht9ga/ALtht9ncUcrpAK9PTQR7Mx3Crh0bcWfhyrInF3Dv05cR
lhJPpjRrnMiAoLiKKSKYcJIxF2HJWkWhZVt6CHPkNF9pxhRnWTuYOqrztPxRX/Znz6LQfBq7u1rj
7kYyzVsBu/M3VTqTHC9fRPymCLPq/ibJ5pEixLgBonRUVhspI6YjFMQFkHDKSq1oLsN9A/JeCpF2
OmYGpe2KECnEycdNQNfilLwKV8bleZMKaYX14qFUT0tenE8YST7/RdCyMKdSn43yQEc9qsZJMwwd
oAuw9VwmEabqGR+wbEHszskPltGhlx+es3obXjNrSLPjfEsCGrT3jVolHhZUdgJNY1pXYUEzmEV/
Z0TfZyqgl4QTnh2lQF9kB9CbtiWis/PyNI+O2M/5BX/9GQR1fL0HS1Hrhbl6l47qf6k6cdJf8RRB
f/KKrNVhbOpH9gyoHgNjnJUf3oqGXG9aM4rstsBVrX6JX32vOKQwKHWyjkxQxXQQTW7e8b7IBu66
m/mV1jtG6XKNhpiZEIuCwpBJNr+uHStDx+WDXtq37HihSeV+qZmlttNUzP5NOj7dTWsQ8cXeD2DX
Xcv+5FH4EHMnJ1UGRK9gBGOxpR+VQ+H5RvyayaoMG8HsUwNpCBLeVSv7FwS83u9r7VF+Ib4GKDGw
r7Ix2teJHTgKJLHfWq/hCpbE3ChDWAs7oqPbsoWwlseSylcZuR2PawKCW2z0sT6SoGQDFaEHthEL
1u/T4DIWG1HS1tVNhpKLsr5Zs96i3oXrjuLPAD9g8qOTVyIFbTKyQCpMCJIm45Aa4XYm1u6e4xI8
BfVDQRqfJMZ6aKFw7FDIyJ+XyfBx7RWy5hLAgkPmP4rRelso/adtU5rpobNDFj21VDQoq+nK1v8N
Vgt1nMS3epX1o+zpcU6S9yZwHfmOxqKWyuD9qTA5mMmLFCYcXHOt1CMO/l6wx/s9rrxv/PxlREmC
DIejfD8pWkAKf0zjdb3YAdSNOd5bx313Bf2+/kbHqQX3lHuvBwmjIwRHPNUfDbCGNzt4ppxVvF3F
fGpyQpMrk+gh9tkrij8RbU0iDpSX2guwh/UhZHXRIv71CkghT3uuqIptK7R/0Rw2a12VUJIoB28G
q5XOofnNjQtjkhJrT3x08hx57zNqM8jHWvImKCKYw2/ZPreg4V+kPoHkJszNd4qFwtu54VOyQB56
8vvMN79JgLa9hRnsUSbA+CSXc9EUWiJaPx0Es3kA7q+XUMjall8/VOf4lk1CFi8lwhozgXallpXk
NnPJpuHbgNTZSmkPv3Qyk8/kH4QnZMCpY3N2S5tWKb2opdzmOTbH+iFQlBFdo5GGUdd8l2BYo8I8
sVcii8E8FP341yLTr1OeH4SN8xTlS5Y0CEveica5I9yzUK9mOurO1z6B0PfknSj1Umksp1qcRvvv
L90Mtju+ahsJTBQBPJj/Y35eqZqte4Y7wSEFHUbGJ2p7mjYK5Z9ug4xDHvQBpS8XRpg8/w9PeKFe
o1W+oFz7XflmYK4a3/qvlBjTU6Athfm3U+GBcQutvELamOE9bIKd10MEWQnFVdZ4v4X7mCSMaQYa
mOzQSbjL3ssCWs06xoxuVYi4/0Ei8z0EqduqMt4kAHejO+fqDEud7s/I6SPCKsg/cN8KfwWbn/EZ
OcS20n4i+MWcy7JPs8mF6FunfO5Umdc+UMI2qaaEZMVJslyeN10vGbKfxs6qnjwy7hQ6K1mVUbWl
q2zciORChsJk8jTm2mi4Tg89b0izqDoiliyvt9l1p/us/JRhH4Tw2UUihqg2CrIWWPip4jLFc2C7
2fH8fPCG8dMEYd7wYxXFdldjAHz5ZZh/jxr23msQenYqNt2SUryxo1Lhx4HVf8ptS15JgD7qTMn5
+mJtzXhsWapJGK252CjgjeCglWdB6eIZ5kG+NbHVfAYCxLFZRQKuhPB4g5PRpv8c2LSScdnuYZaj
LQBdBtPfteg5AyUqCvEHNLLIGdVanltIZksn+cV9HDE3J1QCWC51WS2f6AdPU1zIeRwav454EP0x
9BR3fEz2TB+DoxqJ6ddpRruENAqblNKB1PN7u0ZQZL6TKfxPez9YFSFxRG8uuDlqYFVOC/9SXmK0
m8zc+A2XeOwwoXlBDLhZOtv4uj6c+5yyIABx0M3MMY5DanpXz061Sj4EOSAfzZ1nABfussqxJU4s
eZsNqmnYFoNoLh/iWRY3Rex1kUKukLVBLrwR5kquZUW85DnzAaRad2sf3+4j/0Uzeb4rOQx7OX1l
sXhTBckJ57JmvGSVA7n/j9tcZ1DILsPS2Nj8JIyJuP4j2B0n6DN/+V7cIqKVcGvP1+l2rdxlhD4D
RHa6g1+y03Y3B0l1mOx97lCE20cYUShOA1gLOi5qYFUKdVI7sVhZ//x1RDk6G0F4WWzbNIUdbc7K
aEpukeAeHXd49lyIPP+EbVKQ3HVmFowxYSnfAIZNKPN8OYGKcyQUaABqyO/s8udYU2zTSdg4tlxD
S7GPqkuRnuU7+0jbcQKpr2RBP2p5xPaPl7ZXbET/FOfYce7X4374IKlEY7XNsUX5uM9ycaZhUlzu
cIjLHthGmIrIAakTpIfqXj7oQkCDE2RJW7sw8mPxQkk7k1Rtl3QUdh2Dx/MlEXzcTx0WcnQytfMh
YdcP1T0KZcYn3+R1R9qPqHUAnKzKBkptOzxDOnpJVTe4GX54CDwm/CM0F6cqWqjT7XYHDk+oz5Gq
OYnpH1KqVFMKW1dHhJF3ymxfvskhuJNVvQblpbZ8pPAVwrY409a92WW6rVzGxmlBHT/Gtyi0eenC
IU+dtoh1HJReRvB76QsoWi0+6sd1F/PEFjdaXq8EctAnuDQmQ3xxMUilScFGy7eak5UJPT+6IYID
AmhoGF7xnP9x6f7ykRajLaC0qtjK1EXPBTU9g7mMzYfzF6aCPzj+oblBr6mreQM4fpmzuvZzUArp
CdQDJtMMyhlpx1hAgzPQyjsZL8zCuYJwEFKzPnKd/0DpxRzlAHiFBiuXP6Eb0K8mpXcLz4x2IBQu
N7m+b3HpRQJ8lwooUG7sbgE2YFYv5emh1qARrgS+DO/lXGTQfcsLR/xuHyP+qijTjnDpJnFAtruQ
krzVNidhxQrWiclz+oUAiI73pa2XQEem09eg8rOAnG3YjwMH0gExuxoPtIg/3Lhexib71uW+XeNV
NFWhatf7nnjME2f+3dJyzl4PjBEThWlpJ687m8vimq1sfpJX8fBa/yA2ni1lRXqQh7Hyh61oCnmH
GIVz6yMhdvFdP7b8uHxgL/KT+ktdLMZ5Q/x9RvZwOGrROiONGSjBOZuv14M6tlqW+UN4I5uvTNv7
ybLX1Kh6WXkmERPqStuRAOj5HkfV79b5NLsWAdeZnyxShXv4YQDmyeOPhdv3PiwBiKB9Gn0Kv1el
VoMN806+NKXgvBvGXv+BmUrLH7JQNZ1QBB4k0tdGJY4ypirfhP7rItvG9L5yt08Wm+GczmkBkFJ6
uwyw4wrVgvhz1sQh3cS+iov0fFYQDsyeGb/1JKDBkhCHuVovohNom0I8I7D42iepLBCVLpE2aqld
xN3BnN0QUKZSPOW1pvaSWdZjge43PwSRcZBDb4mPs4MWwBTnCnZ1p6dJqxlUjmWIz5sbGdNeoQyx
cgvBf5NhzN8irMCa8Opp+A75qm2CK3qsvzyemxxRRbAW/1aHnbF5wGlvNigQtY97SR/5JgMlwfUi
wFRx+yhFDmdAr1M3CclJphyo5QEofHisHemzqK4EfeDkFaErBMa+OFWXVCgHMYexT1EXGT9a8uqW
DO0N6oTbZ0FoS9E/qMUXrUfWZkVjcnqEbdHE+GX/y3VdY3ax0+fZFUFxhATsizwAHzNdsrgk0CI7
IDSpFYrt23o/AjfMfqd1GzIUWT0OrDzqnh+7p7LY3LMjPoofgICJtkG/dW3bBXkawQBRdMzY52+/
lj/+WOwByMzXKbk6/79R9LZh9TxUQONjt8ufX+by61MXPTzFAu67h1zp1oKf30WElK9tXmzf5HC5
9m8WNmDUYT0efr+LaOQT5ItyIcSAKcoGpJr+Yjum0dTUSHws6Qh3AFleYTmeJqy5LF4DxTaaHWWN
cslw3pzdlMd0O+APv/MGhPiJhJqELWLOgBwGlWXK8c1CwGD0b+twl18zvIcuy4XUGDLLkYPsiQm4
NFQRSFJJ4lqSVjtya2OkDd2xtthklD/iSk4ZbN3GLk0NTz/eh34eOgVELnTfzOaKZWitehTmnV66
bk2K0sVyABH1vGXeR/7NMkCpAbyGKkAK8VewKkmpiPO6ySolJMvpT+qv8RVWCKRod/5HepDlIwcK
g9G4KQ6fC8uHty6K+8EH4/ZE2eFJbJOv8gVDEJHFKg/lRjT80Q+IJihNac8OkbMUVhN1gXTmC80f
6PVCyOi9Jm3dh6wshkbfVqNyQk/grpdio+uwka6+JfbcR/6OWLPpHlCqhpgC/3JBiX7ucZY4Sbah
l2j+q8n+FaXnimqI2CQyEMOLxTk6yawjoRHycLlS3uaZ2TiOKbJfySRyIFUTSugaYjhyA3PAw79M
Mb9/eQ5qUFWovcpXB0Mv0ZD3ip5aEYCfcBacwrzZvk2i+OnqCXBnuNAvSh5bhrE9gBjc8gRxgFtU
PX7s2/y06PzJYLUD4TrKh4Tkedg3ecnl1rh2sggd0FMLAWXAyqcs4ufK6laiD7noXEAxlxgI4L0J
qHtYHc/yh2WFOqYrwK9QQljQU2DAdKmbXrnxs61jXY8eVQ5xWjhxYP7L4k+XMAEf3Kwr52ftwGmG
0tfiK4jzSgeKJlPKU3ZynlBQRHgQScYXbzJlRCt8kjYk6fMy9WYviBv8VGbTyID4DpXAB0CENqCD
SlykzliM58UdvOoQMlqgIzCnqkoEUaEOZAn0T98BdUWdGzSFIe+26eNvijSFJAQcPJaPVa6a90k5
lRMpBs1dkt8srGsDcdw48u3/PEOKGS7GpJyGdp407C9M3hKm4zpvng2StxF9r7d8+3axGqepgloS
jhMGhvs4ohuwiFU2k8NLtePavJSwfEqbtv5JqZ1BZ1fyzmeUfw6wyFSjjkkb1WsMSdfDO2w7Sdbe
1Hm+nbsG0Xz36LzcM91Jb0K6N5VtAfLXiA3366ui89FaicBUj8gPUFpTo6qd00qiaCNi/D1iCDod
eRCFQ4ZHL8cMNOyUT5UCCDh28HSWgeaYjJ9lNHedPrYFP4fSaWr+WeqHILzc2fWb9eTsc1Ldk+JI
bATXiwYjEDZ3rNaYzsdD7FN/ZlJ5NBa3ihdCTUWfXISUe6V8J03+RqBpgUbHfdfWDLWn3MyG1IlV
433BxxL5XeGyrfJILsrQb4BBvAj7GND7A8RHVagqlmhoLn87euLbS+VQICK+fansEzH9zsGZLxNY
bGUMNDZR1uP78ORkNbccPjIAu2Cog09coEN1IMGsXglC/vG5CLqmRtsgQUIyg0fLXeNT/qGvSpL7
yq6/TtIvQyk1M1SGCfpFvj5mYLzG/6b3XKLIw/yXQOdMHy38YYw5kV2L6GX4nKu6NZM2MX9VWkYg
gbMeOu/jo1tmmAiRDZqoTtmkB3wr19Z9Nf85V1U6E0bsOTtAq03+hLtbOOhCOO0B0Zt1wzM08orJ
IFZtcdUwBd+rqx6zrtZ+FRJRLVO85xWwinYgv0M9FiyziW57rV9TwUrgQTauWZMK5DrBSD9p6ZYx
HELWkDCN76Ygu4ffNcQqC11wDI8GvRwd8u24J4stOlyZLyj1bfzOznoqkSo+RN58dUzNhKFvFUd8
5BKYeb3TcvFYlW6+uiyMyBQm2BzUNgOTj9njZtyyUUR8gp6UR3k9Hd5bFTX6VlHc8CgRFWoGTfpN
cAqg+SDD611xkZ3VD5DBRv4F92w6mAgIsAMPlQL1VtqleCgSPfqIn+2jF2EhSN+K0ZSyA3QrSg2F
3n2/JCiVzpmx3Zaqk4mCoXBIbvy4Qi+0N7adFDFxbzTEYV05QB736M8ikEta6W5RfLRStl/OC2az
I0c6kWNIIHESULxjzzyuU7hqhghudPTkTWus1JDNQDkTRrYvMPCB9Gwz1n9wr4OL5pJK9+6J1HU4
yLlznp3xa0RkvPX1RnbqZKXG4sSFgqHrSKm7un8wyXrhUEYPilMB+H7JXW7B3768janKmqheV6/N
h1DXh5JkBeQk/Na4PaZmFmqr+zrlIDkkh6DkcPpssLWC5oQ1EAhM3KAj9Kh6RI8b46MJedKiEglv
j+a6ni623s+iRYltF+1K9EOrRcPPEI2WRq+z+V5cZDsO2vjigdpC6+tldYTUfDi+4D1QuutKszgI
03gpxb0Pgm3SrGv39Qdi7OYJnW/dZSNLsRJBogoqeWq3y/LFH2GJfrvKhfQrVXv4dUpqmPu0fy9e
4w53vYfFDB5qSw9C3eAwrcnfXFK+hEXkk/el7mlVYyB8Z1UVxQeCG4vxDPoAYXITdZterl/j63wq
Ui8nqZ6tBhk8807ZGNjHAshV99bfJbU17PWP8l6o0N5uSCOeTIZnC+a+V3kHKddBUiXs9C4ZzmLI
biQtiKpBATrqkmJlBhFg911lR/Sls9CwCgmueJV36HcUm1girSwXCvmcAznBJZMWQUhLJZP3jJsw
FtWlJTysiqUM+W7D6pxcCTET2zLaEUpKKZkLI2wYGvakHOoxu/VbxPcRTzGg2shxt5sz4E8GoNMz
xogcgulPNe+W26p1K/1L8CpOTwhxiXoZE1f9NzygMjx0s+9UhjRg6uGqFH+RghLINQosQ2dq90VX
h/lga2XyMxSZUFsTxoNKBtTqi3iOl/M1KwONR14/k0HdVGQ41GVc+KrDMx3w0tMDlKx/mr6tm9eA
WKZE5g/Z56zqgh/JOI6k1VKq2Xve99CwSimB+6v1hjXgnaTqaBVibo7BPE2sh+OVjgwK7/kBCRMr
Ln8i3XXrkwr6i9Y7Ib4b089qphLsAlwif/UEEzbUXfKdrjIwcbIuxulRnmYknggRhTj4cedDZVwL
yJlQee4x3UAWejfCYoSV2e8afribeB4HR97PxPo5V/MUmmAHLimlQjnL5otlkgrZJgwrJar8JL0U
Re0ZtFqszDnp0+I4uoHtwT5IykEx0DYPNU74+geIYy3wW259o7NyC5JpfyI1NSkMqgd8VsVKd3Yf
eRrG6B597H5Te7XnytfERpjVA9/IVYzNgf7EgbjdyWxZbNxRRnhdY9SJz4cKhQ7y6tQ7lZxLrOlA
2qy1ji9r5NIhCZX8a+jk+gIjvOC1fv44wpC6xlwokGEF7vqH3xPjexabIp+QEYE65ghV8eWn2xiN
4ORiAWpE2Blf6MWKRcp8jIlDib459z5YrIYPqxpBtSDLEB6Cmy97WPd72Be8Co7RVXHCx1blJZjU
3X8o23Hn3TXJfgsueZtHZmWUEaVg4HVjo5qUfegEMJ13PdwOnlbHPZnXJ3J0Uf37wHCaa/aMVjSF
jkGuVbhA/q1XcHdO1LNnRN+G9H2JsYQsCVuwiyeWndHcmPG2NNxhKfpU2RmSDRgZEK13ES1Q+BJM
gQ0DLHmZzMfKJtgbQHMbhbbOvSFJOJuaAYZi21iMaSjN0I43rE2F8ftywSMkiudlrRvaNi+buL0p
vdwwm6kCnTitYKlYiVyzlcpZ0bSgjy1RhUDx6LyTQW3rP/9XCnWqZBdbPSyrOykcriTOxS4z4Mkf
2EmgZ4YAcy8WdqSCp0wxKGynd5Rwi/Eb+FIIOVeUVN1QiMyhrjnpXO4/vdg+dJE/9riXODHkETu0
nKDY9+Gafp0/yMZL0VQb5jbxwkzFW7dewsC1vniSZ2F3KGLmDg+JZ4Tpan6z1LaIjVMxl6eWlXVp
fPrAT7AMeCbsiOEH84cvHkbBSJuNKfOlxk36KhKrpveg6JROBPZIihzwQJ+PKFrZcVapFXFJXG+l
gPmpAHex89ctRb2xeqXjSros2wovlr47+CXN8wQIk8tmWYmoekdh+7ddYxuvrIli9KFdT6czRUXa
dviXMjM39tr73ZG7D07tRKOk18lfdZJ8CRWU3atOyvMISPy7LVxDAOrxdv/zx4TZ+wDyxSOalyQ2
btGQd2zAP0W2d4VtL8LLD8ivYJxJRPBmJuDXryDrLKHFvsNVN/g+/zkpr6M/GaqG1JSsZbYcMN+Q
wTwTB5Zdd3NMucNr9AQTzbE0fp32Cz3W/3UenMfmQaLP4/Ki3tAhad7lwax3LKgOhDxfOe+U0bao
w/XXleWKrkkT6up170PTwr28fFXyYXcAQwDLU95b5xUZVK2KfxWoaIXIg2sKxybFsEP1Vq4D5QmF
k64E1cOMg3P2vWiHz48e8gKQUVu7A0RJZGGKzFWZABumI/xDhMVixxF3ig8ALncogBtooMhjHXd3
ECfGlYMwFdRAlb71uu745Y/wbq+P9j66+Caz7yd5j4aMO5VwAAKwDsZDvmebu2m7TYEp3knwVgoh
gkVi8cWakF3ieQOF38tgghXkz4Fyytwjhr3fZk51CmXtCZLP5OWJ1KwPFGFal3tehPy7Qm+cnh30
UlvAHtI2dZKzr2W1RYMfg8XYBgQHF8GxKdPwYi5J8h9ExG/lLji6QvI1hYlDeV0tcBDkUuolK8uj
DTDyyXKMw9yv0lPq7mjDTJFoYbodUore8HdsCRu30dfBxmSr/2ZLasar4o2lukcqo2/592/lBa0A
/+5Ri/QpARs/FpnAQDXEMpnwA7EWw7NHxTqRL+LlzAVQy5Fy4xQBAbeADQJuKW8n9U72vk/6v/ow
rtvydTbUq2OAZ/1JWv6UrVk3w31x6yNAs5N44TLCvJSUS87VOoWEUs/MHHz7KX1Is33gMQJu0JT5
xcHH5sTif53tSJkPhWjyEb17c9F5SYN4DHMldEOK9wCzTtkrINoPLy15nQBU1A0N31TSXPDT4pQB
6DfgZV42XRu4/UB85VrSawBaFUHJITgdYAuYsk0ddEy8G+PqYAlQCa6HRZeCyxuyOt6RLiQIe1t5
i2x1pX+ucNg4QcdN+Aaq3HuyfQzsUMA0eBh+DIGPVaUbURT0kIEnQuE8PuIuFCioOUYog6LSJV2C
oOjTGs23LvZN8dsDByb2sIWVO6UOZSLo7lisB0Dhuj5nJGAR7qrMGmUI8obuZto/I2TTsfZTiFCF
WCKggOEiBA649PyIMlvqDp1IvulX3f3gTfC5d7vAKLahYHEpuPJVbgsUCgLScjOBjgkp1gKDpy6u
K3pqVF041M5RCNPQMzya0gWXGiqI9AfAy/e+lg7RKNhHHkYDMewXdKLYeeFsjG07sQF5hhJeGsPE
pwK55LQe8TFlvCnogPtu2rQiHuyUN5lHut3rxQw+40T767dOXGS6M2LGr/gqyb2k9hqY4UC/Tu+V
puWTrj1Qs9AeQ2zaRIauE4uN5eh/tUQw3cpozFj1GAFlwOx4AcBMMchlIYD+dQ/DJzFDUXyzkKqJ
dJ0eVu9Mglft11uQ5V17ZSJsENRGukoG5OGxQGaFPYPRMJGEdQZncD2ZQdq3g62a/K216vs7FTeR
4nL0HIfa4Ul31t1JjpNRT2oqcTTF7XqFGJPG0sv7NnHDo9U2Cn2ReUNz/ymyZgmCWgmpPB7bh0UM
/H4XxPNHz3fePIePLK4UtE2x7LWKY0eILivhMEbKK+O89LcCvaXnudJw3/lnYVlVrzAx0sS7j3cw
m1wYXR4mqxUg895/dXeUbirxaOTsXG4ztVOpjBpokPqrE6atQwiJOAdg4jVmqIQL9V2u0ehZ/2yh
lKkxB2Bj8stkal8L/YoStX3e6zraQ0UNe5ASt6uXebDZi9GJAsODIi1TFLUdo0QDeG+wg7phkn6c
DDMGSTJn6QXqYn94rbShIcaKwdle929CZ4KpZZiDhknnvcWdqOi9VwwLAGTa91dSC7VvQ0+16RUl
+qON3GOoXGKs7SCKz7Ig+tDQfjjsUOjdS43zxHtSMgMfHvmkpYGrMg7xKXJm6JxfCu6ddTDzVlgD
07Km4MAVXftvcZ0k7FH3dD2Amzym+C5l5Cj4X21BWFFwHomyznl3dDXyRK2/jsNV3Yq4A69G7DT1
9rqoqIsRAytnZ4QSwC9Rl5NVjXbEbURT1lrfC0TIGvFeT2HiMcffCptt0qAHxfgO1SUhnhycSg1t
uifTgS0y0wU15Zt7jDouoG0p6fhzbLtqlY79EXNGmd1LAhymSV+03JLVxF+eWM65pfNGlUEV0E2v
VRKo5iTIWC4ngwtY1ZlSA8iwebBxedWdc2g1MI48MuyRVVbRpgKSNcIN9E9OptfS0byckl140Lx1
2AL9PiQpm3LkC+yBqdMxpK889F15iM4g9hAoy+0g1AJZO05cms372JXoXZOuz1n7AyYL/6FaJ+lS
PwdzPznKm4EkWhoUFuHsPjQ+OySKHQuqpOf7J92gGjO3AkjF5sCvitUyLxsgtg5y4XtfCmcn1Mkf
naA6TUMc1kmAr7TcIk8ROJ/Dzw588sdPsYtGUhMQ33K5dbsSou/d8CODXOOokAOLY8FJyTcQp0vs
ArBekHYs8hoXu9gJ5A507tpU5vv6YWuaeiL5OB7Jxs6NuUyUB6Vekp7eN4NhXKOse7ado9vS5NVM
Ljvo3ZHCji77p48QOzCFlr4XlPeptdVY52jvvNE3MMTDQDnYmHiVsd1bDmRGQmQf7tFapQOskZDw
JQxTZzkY/vTx2FiITYkgbI/qnWkPQS2x0C4WX/RVibArevAC2q41tO/i1Zl73tf9ddbsHxO/OXSX
k8SnDQlbx8yfZSUd0qpLYyhySPIckJPpuagwOButnBEddcJukSbPt3AR/dmshikt3sJ0Su5SkG3V
+ovrKOm++vrl+8px9CRLxbiFjU6J2xr8tOF9q/InLD/BJJIi3okfdkfd5Th234/wcKjCvd6NKZ9e
JP7Sp5QaOwxrxtFuOgifIDlW9C+WAEiBfqsnSRGA4qUqAPaK3F/mR7onrqtpnDMIq6jJmuz6jVBS
Tzp1rlNMBrUm/sm5akLkWxEDfAZ6EeHb3+rc6cItgwsE1M5gT4zUnkHoA+pJja2E54+FcHRhv2CS
x+srPtoLp4hntRmM0GvUxhy9D3twKTp0Ya2e7Ih89jMVsi0w53DBwhlY1EBNl4HW5bpnN2VlAPKD
opv9lGeBmN7C65jxyTiGVGtqrg5VyNeaGfWJ32q8k3oik90VvmED4ej4S1+lqrr9rCnrMOs2+BUu
h+yhEBf0mD+wHgPuGLJuujJTVhdqoG9RDRfu3n6hnWvI6RsUcrSm24jVBaxDjreBUY8rT3SgH/d0
c247gWjDs5uNWfWR/LWSXWPOqQTaO7apDjlEZNkbtyIFqZ5cmAE0gFKdWsX+mx95KTXpHd2RVlWy
gXhrJbWFJ2tswxsOmvDbM3uB0NBUpnuo4Ik3fno/Yx5PnmR46pkAyY4X4Eu4tAPxy+dADaKkJJ56
DVbUWQFjElcQo3Z5wdI49N9UTMLmwGju762yQun06o6QN1JV2mnCikWkYU430rdxRSsWufLNu9wa
juoel7hXQYtbis1AIkJP9qYSIieM+Jfehv6Ak5bfcqWEQP4L6MQE2qUn96Me2mH1jUHN3ylyZW7x
4K2XFq1DGxRexZmQ9ZoD2i+fsoKJPtMC6jIYWuaWSbjOYahvrZk5y2Wrk1HQlEFYBLB0IEIvAC4T
E2nwpJm3wZ8+vxeWDqt6/zSDTdUbRzxK3EMiI/k3dCA6L5B7a6DKmLwZhCMR9uKqMLj/m7VBIz3M
B9EClek06IC9vFNHDzaFh/UOOkx6hV+KqRDFsHEe89pUoE8qoQ2Jh4c1KCkZX9IPfibIca9xgCBB
WssMuPD8Qy9gfi6H/445ItG9W0cACrZ8LslSPYezADdN5mmwGXgfp2QDzk3qqYGOi7VTJXSqS5UA
LqOgjhX5wmxjNAoMUvnCCxumhpetithCwZf0xyi4gp49r8j7CUkdRdVPOsTSytUa8+jDu1nqIGkp
U55P3tOFCWV7GERj4gwarRN4Z40YQ6czVLj0c1htVuNx4XJsQPv5k8KLgZyVg9FJWENufoteNU1i
cAFTDb5eOX/uoekFg4hD9qYowbzws8p4q7rIZkMYZEqZWWeUe/ujCSiLQ38kgeojz6u6VUaLLOaZ
I7HRnrpgP5xDrcDOzltLGVSfVVpDNV8UNpdZHPSntVVCGznLvPVpN4GSCBNjaG2CiGJhpSTlsFwl
IiaW2QzKYaOSDiuP08GFPXSM6IQjpAYFSag8q7IO8JEktEwP4wCZAbKbopCILDO1UvhvOC7Jv7Kt
rPPHpl5FEzzfQl9T6vDM1fL9Sb+4Qbcy2fstYN/K1KXSMPLYP9T7VU02lHOMIzR3nLz7KXSaVSH8
JxyREvDjdEO0/UiQyV1N6+zZtZrgp8MWkjkupNQ4NcsnaLxp5ufQ0kL+X7amWPDD2zaZfhCL3yie
CLMA0FxgAT0RpuSluRudiU6zH68vy+QYq6V0JoCN+neH6wMURHqqfVLMM8ZuwJtzCZQp1YC99GN/
GF6OKbHn2MjR3WY1P+uELxbySM/IZEhB1jjH1WV6YvRZq+7BfNzUkNZVYG8ct5L3ttDIommdJDiu
zbWM9gHwpW7oHxrNMLr+SW6tL8oq7WF9xnSXWUGSA+i/Xe4UIuu+x/vThpdLWybe4gegt/NJF7mC
oL0/nLzHMtNmHusv9JyAQ6PRTxPIEa12vTgZ+JP3xW6BKT1qBrhpUFEXKjF58+72RmqbNcXdloDT
JTxpPoYA/DHFvaP/VA+KnhNsMpvs8LxeBnWMkBq921AEHNwPeNFnoigzGzxhV8L5yujWaYwzCVmY
/tKIopHMek5yM0DFw6LwP0lQVhQTweynTiPBIUngwhJxNHcjvUxCiPbY02CfLKdLiC85HGZJZh63
B5gjpzyxkdo5+tQYD1alQxmiEBp5puoGfgyRw+AGZaxgCd5JAI1RLirvyqP/zPvnMur7t0lVRPEm
7ilIxVsnWuLx6w7bwehaTqkM74/OBIKhAsuW0cG+T+JiZb1thCUD3WEnuTMiUqXUHd+G0puR031V
cQU8rLmf/PEq/nReTbPvmCtj1syR/JACVy3xHYuGhTNSplQ0rKpBjnWFQkuUwalkhobmyKWK8U27
j9W7DV/7Fpe5k4M50OKb9RaeFdla7xpb3nB414etp+W4HTUO+rQHi6FkZvgBpc0zXUuk/AmRhLBm
Ikgfkkv8fJkFNf6uCom/22634aaJWmrqt6FcBxZ890MHGHwHGS4LBW8xl5OjsZrhBppO0/v2Zhb0
ev2/WCvC4aPK03oZzUFCjnXEIDKM+ykmyil09bVPTNnqJsKxsUy9c3d0HtTc15zsESMvryXpiTvx
b9rLjvIdZOTR4XDAP/ZJIlPt9yBLcm0e3jD5E+9n1Qr+fReWe2/bMYZ058bwZK9YHlYG/bvr5Bga
OuMoKVu1gmlav56aDSNvmYSr5mKD+LnftGY0G0ndIB+ApNnGvv6NqU71LCvVVXZ3B27g24XpicVU
uBT8jcJCsSXwmiubGbOERE65/wuCQtFMH6bbNKkw8PuUE5PgH+UVlIgDK+nOrkOSavZhEnnkW48K
231XLS1JA76SvBW5gqgTC4VoMfdkS2/9FbcJQn0xBu8QsnxQujvixeGFqY5Vk/bqxSeGdW0J6dnu
58yV0+p+qYpyuUnxT7ksIvbb0AhMSTqF7JN9JfMXJ8ikGca43VSLmHPx3yDI4uujRxUGAbaxdPpZ
FRXyGludpLG8cIVR5ZSKGj+c0/Uhd/56xqPGXGntCd5Awp77HZPvrFbrfiVjniFM2Srq+w8SgUYg
QbvJ/KKlYe+dMM+H+7wjWD5TSIxsYNjegFw+V1n6EHtidEbvvac0tM0r3iNNXkyDl/uieyuuTdbZ
KDOkVlAGuR28aZdlhuIt3TfaAMDLiPOJYtnKSiLPDHS0xl/nZgf1fn+ALpxBK+QZcB3fd+WS7bXf
KS5p7x2D36RaRpwdHRpCYrHvXK//6zfXzfzu0PDbfPPrOyZgJy5FayOiWB+brSJxLcGcKDjLMreq
101bRY7lwIScei62qkzb/xIEoNmP8saBaYiEtYgiCZYjl7rwGRy0HzVJp5YuG0pn4c5xVGK3uw+k
VHi6oEocRGSzU0bfT8Arbs5vci+ddywd/3S7c7pmQKG997t6W/4lVpMcQiBeQhi/Bg5J0a7LWwTY
OwJnjwIMIgBU4wR+kHhVTlRRg78s1DdKplwpbYp/fIIZe2l7mPVZJ9evpnq/atYO46v02k2udkPJ
PAaiB0KZi5GgCwr8XXHaPs4sXggS9zpLwozMNJZjfVUBPKFubvpAlF4lV+NBrx1lN0GoBIq0JEAi
cRe9Tjpqkof7P7Um6qAU0B259M2fx/eZxp51RnE9yMsw0sM8vaINcgk5mX9OeGmYnlfcgcPfo/Wb
w33UHm5jTQCH5x2dRut/QhIb1M3/LfMb6MXqRGlKXukXWNFKv0ZVLax7BB1IkIC/43+zgF7w4iT1
dtOEHi/6gnlEOJkSCUizCjMWgxYzskPe+sNQQ8o7UuHZIMLL+dC0BHgtOgL8ViQ9HXPvmS8EUUQq
2rfOAXhAZghuvs6do6N3pkl6AJMGfj4vTQ1gwDEjNSaCp0D1V63cNfcYqtzhlT5aXgNa7A6yLiqn
lH7JpDpf3UPBVSYd0NN4vIOZRpnry6hfcc/+OquNFuv6SPBbcHIPHTYaTXMVQSmMsjYy2JpvpGjV
LSxqjOuKqJL+oFiTCL7h2KzXDrZ0f8QbIA+X8wQe5IeMRxHmASjww8/e1LxH84DrhGf7Mf/oMo9y
reY40ms1tRlhG0Eg5gt9ad/PALeGXeLiqG1P35CSe+QqlI4YaOqs7ccFy8S8LTo/lJfFPiWo82mI
qOQB/k8SME18Aypt54+8SCE+M7AJVec7luA8NFr2MRUFJbJ5ZG6oM3WxPoAFKsDd4VG/zIHB0zgL
Y6lU7PG+HPsEalT/dEWMApjUp+quSb8fvHl0Y1NiSkYgJA5uCxSxylxevjAgh50e87ANMGoG/4b8
B96g1qT88J/7AW49025UB7YJFakuhuONXFMSuBmdxBouZxe4D2y+wo5F5oEOQRPAK4VJAxmA84a0
p0JDsH5eiTSAtBHpBu9xNrd8mZih8pvvWTo/9pHDMKkpwVVEvjNhk3ypwoHGhF3m91S15uILOpl8
8WzH2he9hgNx4RafUOh+9Lm7fSkkpnqkNROzQzUVYHqkMf4sOSTFQrgXkM7nnuc6YKA+a4ZDvb/T
upDICvqa6CWFNGkpXIDpcjve0alOa7yO5wadX92rXVwcNBqMweebPI1WH7HOEF5QwkyNmJtWknHI
7KCCPw1gkWIUJg11SbwjNmj8LXIjuW1+fF9MVJVyvyLvSfS00MRlFA45gF6klSV1dISmlxjPtnK/
XDFFzAeICPUWXztU7+Ss3Lsv8fK8VUUaEO9cXoTqSEiSoJwpiBSwUI+8l4XXdAuQPAMrNrxSrwRk
gVcrUjh1PE0dGqLsSGmIP/hWE0zDGnMs0Ms9mQw81Bw8eipcRLUN4t/jlbCPUFP7cgWuYIRDB7BY
pSegtkFa2RYrVRhZG9inyNShdOeimBtSW/1ONniu/cjxlMjQsFVEdvkDou28GZTCk7HtcMx90GTR
prQzeANLvV59muwbatYWs8JObsngf/vCoPmBfe5BeG0TaPN68OwDY4oFAQNvfMY8lNB854MPJhR8
A5hxx6BiffgW0rwhAaNZi1YA2MowxbbfQu5tKEU6KHLzk433C9ewfGNNV1KkKro6dGncR/e1bQH1
DlX9YsCiPlDIX0+hRXqWS7F2k1HhjwL7PrY+wCP6SgtxArCjIdukSK1kjC8Wg3XMJWqeiI8Jj7hV
W3+8uuNpzPLQKi91jPyVFRjJQzSyLl4GBhWtEr2nJjEXyTgTcCy+x1MuHMLuYoFu2fQCyVnmLqOQ
wgIQYcvRWLOM62hP9BeMwtDNpS6DMDtNBWzZtLGadi2Bo9RT5RcR/IPvloVVMpRD7PhhzHy6klZ/
FLyMl/IyO7Sd98XA5MrfYVu+/EpfkVZh6af6tqVJQNHOidC/DNFkzQO4U9vH13HHEu7c6k71I1y/
hwVue+sZ7rDVx/AMFmueFpSsAuG/1VILn9qSTZofYGPVm+CP7lfioXSyTkH9EkqZCWJ2FVbJ2MDU
tBBTfEeXVRwoVsdz2608JPdbJ+2OGvWu0sIVX4hylTHwpN9AnwoUoZcvKOT2QNOoKM4eHyYhjAW7
oKygwK/T7hNMm+h7unePZLiur4WZqPWkD2mvOr3xT1AVqVkNCz+KUf2N6lXK1wr2WTfcBbFAGSIq
q8ulUAxUkZKaFJK2CTz+ujwnhNX8fFQ1Zfavudev2zBki5qygW2Frncyq/g5qR+2LmovXNFRFQX5
NvOVo0ClbHP4H5yv70Kn4QUTXU3VacMuvc4tx/lC5cvmiilF30vjr4KQtOHo/M59N9CyGFkADVSi
DqYNAMzyIq44OIBGyQU1kOIPTlI1WAm4ly+oWOUF8niaGS5PAlritVXr8EEn/P0WjMIpe8ikkjoC
HUywgJlhTtFpHQ8r0Y3f3ynQsRxKSNR9MkG/wHkJlcwiSvIlvlu/A4/Ae1Dd6yFvYoANs9slNQtH
FHnuhTchmF35pzUGX18PKueGP8SLlwL8wVRl9IqGQumCJd+o9n9a/LJwnsITdSFSyxUKRBlU+GAK
mQPfuplSYxSWUU+JTviOgf8WmBNUvpLysbSGpMHDPMeFRNP0B0c4Ic9ugP/oLrLrzclqcM3mg57x
rm2MqJBg37BAOiODTg9bvT/Vte+1AnInGAL3Hy2hXMC07ibQ/TVRdVM4DnZUwmWIzczVUnKL2gSM
v4aJet+Enxt6rkj4D5mqYs8dFDtOe3543+6B5vFT1//luIh1rTv6Y2tALxYJ3f+kVSZkKtalDY8T
7sdt0N+q0PNvWTyP+lYKqGsY8ikZFZsEw0yI4hg+VBIQWI3yyd4s/JHMrvOXcHZLr0TChcD2uozE
N4r9LW5j9nHpAcrTSTaI78+Lh8dUkd/USkDM6J8ZHYB34dcfyGkWyo0WEr9Fca7pW9feZxEnIOCV
vBlRw1mkk3jN52Iij0klP3MoEC5jkppObpXb1Dbd4Decy5V6Bb+VWHhoPFjKhE2nYhiRCO+HjX55
0g1qUPGYRWOO1lOLPZZwhATZwvseL8j7r0wCE3LC9ekKREorZx7hmw5/e0raAFiuFSrd6R2IQxWM
V8Z6xFB/5LyW08i20A/8GZzMi4pD64idjCYQncXV/WncSzD6MLcdia9SOCT1NdLJH8mBMII786zA
xK2eXZN+ciUgCqpapdyIrDyWUqUw+EJWVPkqjHdvIqqhhDodyHKBL7uViVybevZwBje1ym95x9Eq
vv2A9FwYU251u6jtErrB2FGo9LNjcDL4dNfKfeR1sCZs3Ms33v4XZF6ZnNXaUDjQejNVvnlUOS2d
TPW7JurAYMvC6O6wZsmkE+i3xas2F0SMaE42WOzpSlfDXTK3e9ID/7Vxsx44VdSZoqWGjzLObAAz
jaPwEpjEe10n2KzoJWVRz/TYnnUBAp+1Yflq5KYdTBcVh1aVCDVD5K1bLZuVtazZjrV5iI9O6w1U
JUJLePMyKH52bTU/kg1UfHKHlrZhw4f86y5AtH2n82pv1AJjW0i3koj4jD1KB8kqhuAoHfCWdp1X
RIGRIVbwtlrdq2/TCfWTuGDW3FQAc05WO2vfgCox4BCb2srTTKSyWfFSL3nGovHejrlXv0KMP2YG
SPiTtVwOC/XbO+z4wGyqHr5uEH5XUn8S9yZPP09ynBVqLUv0SlogQAnChnb8JIXw9SzLz+RAge1Y
x/7jLC0TWvGiAa3sJZdfSLhdEq3YyR7Vxu90Zdy5YPkD7EtxxfsOtb4nsQ8ktyiJG2Zy60XQJw32
by/nFSZiT8EiV43JhFd1ujHUg3Bv1UrskrWK1cSB0KyBZHsXIY94o+lUQ1T/VOsGFmVddyaiqk5w
4CAEmE0zGllEO4TWGpZv+JUfSr21AhKzLRA5TTi1Eu4B/zFO2hBNTVJI9zMo6rEUvbMfuOUS6FVr
PBxrkMFXUu1Y30iawqboVXwBWqqU5sTkLCWXLxXf0perJrrLUaMjGqwrXYgLepQcp8MgE9TYq9tO
x9jdhmQUkWQrkxtaMgRhqROTSLrJW2bfvyp88FC95FEKfHli+4u8fK58lyDR2aHfqdXdRiXIwlkv
T6I99vzPSJqe4W1Lk94Qlo8PcISGYTdr44Ts/EZSV3xBCwYF7IPAS7R+Pp2EWfJBu1Sb/hVvcw2E
qcgVMvNQuPadRQ7+SjOPMPXDzHj9YYd9hk2uHLVq/CA24WjTDib7DdegomHWJKedDp2yoqt8X9Qx
OJD6+y2CrNk87sJQxiU/FEACOpBOSV5IAlKICuI6YkH5pWnVCYMV7jx1Dq16t2P0fTc3eRO49s2C
M7FMOuyQBpNWuXl5E/VeUPGRzOpEdOS+bp4jGuxGiMdDVgH/5R7/Y6tIz86+V82NLmbS5x/eAxtv
xmIvHzolwIm1tsf/jch7Puis6XXDiutfAVojgmlUJNwU0HifXj8QIpIzBP/YzKajfbXRKA107z04
/jti5cJTkGDkEKzEar9qnPYjN/crgtPXh9Q6jp6ek5eYop56tO1gQia/3W2OVgmZeaIFOoiqxDaM
i7IwpxCLnU+9LIwDzsuZhesmT2nr2wnWdggeZqLdP8xLvONaPufpUlxkdSWoTpYmy9BqDTfFJ+MI
ijJ0Vo7DNIavYkpNVULV6Vp86TqP0vzll4O13nugEmgHuYiCXU7PRPUOshDxB8UbZRA83aEAh6QD
l6wGmnflYjhBRyVta0+pFkppc8alrl+xCzi7g9+yg3JBjihm5h851eBdti3RRROMjH7bZQhX4IAa
9e2pmFtmC8ODEknSK1/ucFy8LvavndH92pp7UQcnx5BTd4TgLNbIAKvVry36124E0WGSn2xJcZEC
R1DjAFcNw3xJTSZJ1+cO1lEXO2Wxgd3Uq71fhTGIaQZcdwWUQtYZgfymDSgkXTLi0QGGTmGl7W+2
wIyuwCdivvsONZsEZbX2r5Ktwl64K4IqJ447Hu6SJpD08DiXmGZ5pGwRRekkVSQk3WQXBsrMMrrB
d3rheAivEXrfz4KZB8btberGt9UbBzT/gOfUrjyuQPBLg157u3fAezE6ISXdUmRygGzoC3F2gvvy
9ksK5wAD5YxtKiUi+cC4r084K+g2dg7ZhcD4U90fFpOd9Qwb226eAXoW4KtSoZa9ui2xyQIImtDt
urViJZqqQlFkc1TeaHNd5vLIoKRg1OOMS6Xs/l0qvhatisc3NYGg8Tuu99k71ugXidaxrgjW54DP
H35bLBGWyXs0VFjh5QeaO5fnbcQMB0hnvCRgwRtUnhB+VG+9G3SyKD3tHC6gTeC9jmh3dlLeVH0R
X0mZ/NEyOEC91raEyb5J+W9DHPLo0vM/YFvkT8B2Q+gukOY/9W+bmYKisU57/gcIILKeBhpZbQKR
RAcV3fGpvg++5bZ0F5odUWf4WPW7YlatAx1gs+vYYlKYAcC08I5D4bfZ6UbmFu0dbBs736jbdtmG
RinyUg9N1/nfrGbsQ9uQ+OFhg4q87EcE4lUCYeX5UpNPu1w7SZYKH3LlT43COEFzrtLzGwdsKhXp
SnAxZKqQeE8zzK5mnYSPiqMzLwaMUJq1jwDcTbY5OGBxKqUmu107wHZl3tdAE2C0QdzD2oM7O7UG
Gem15eEUlC0EzcYK4Wf6YXE/mGVO5mxDIoLr09AlPQYoLLFPVBZfuu7wfR4Cvwr6efPpx8RcpObt
vDZE1Lz+jitukWfpK/kqWFZ97eHhZQXBzhTzfZPNuD3yQrQu3INwTAmDCd/R6Bh0RLr7yEg6PAuf
cDDYCxQhb8rSXsKIs4T0+z867Rg+RpGbltxSOgnHDyKSPjnfqRecQdN5dVsAuDhNfCQ8TV+2XaiT
BjjfRV7h75obo3AwMq4Dr7vvve6nIVKYtUz3g4yq3xsWqhHj0mAQtHTk0NYkpYMQ19LzrT22dnGa
HglN1OyBy1zNM3HktbH0ju5bvhRpUHxilhdhgJA8dOpmcfwxrlimPQk5aRXDmooNHVGCwY/5Hove
+C9KtMxESJMc/jRAJ07WWvOgs1QRHf+eITZLaPeOAf72KNHG6E71S5zNFmlm80ZTpoykcAVD795h
7P+xsYgNSV3PQaH/Se/xLiGfsgUf1//6Nb/tRw1bZu3ue8CaCOqa6j2nypAm64vhJqtwM1uATqFq
vsV3I7quKKNwJmi/R7pyfAP83iS394ZPRB7KNn7OCca2f9+5zYZMJBURGzJea82VVDeAPWEs9JSr
SKz2w7IBhNusZFdng8jNILR1nyNjnLa6/qX1bZ0kndKjJINwTvlhYeysTHYmn2MXFQkXghcM5wLR
vnPNyY951BPw11hF00pvNwaM7SplIUJ0kr9dt+TuLgv9L6LWPAOrstTi/pQqE//v9f/1nksMWFzP
hTYf88D6FZ3Yp2W453sB4k8Nq47EHXeDpU0Vc19vhaElIrTWxSlqhheCEcRxZglOjVSJkf/RjZJf
lAn4vqiSclQ80C/0VrQ3w7n6DiZdNfgNRF1piDaM0sR6cQyIgDoG/TjzPE+0GmiE+jXcmC7X72Qs
pYQybWcyVSZ+T6UizPO0sLQOaQRUdH+7bOyiXfZ6bUGr9xqeSKfiFij9OTUu9aZuzSLbvNbcwpYG
GfKEQMdCLIzm1DDQuwdh1O9uzx1+wMcV2dtmi6hkyXGlh0NG6AfSlRx/r2oiJhtgXy2z7rxFIOTl
m2as8N2RcSzUYNiNr7BhFcrf1S8Q/nnI0pi6HuaC+9mfic1AaLcbWIR8f3A7J4s7qnPOilPXGgUc
DeswZfD5784DDYp/id/f6tdSwseMihVSrRgOa7ILs20G0QkcNpxUuXB5s7R/bS8nOlSoAuIyLb+Y
ElFLhxQvAE6uqpqVgdujQb3Jd/6iJhpCk1M150e4B5npXtsMb/4qZxxCLzCXC31z/WnX3qtPm/NW
1u4NRPeiGRhY3p0guJPKmLsrHYiNXPoWHtylEP++ff13cXzGFK7TAtYgu++Vu2ERB3713XVup3vy
JPVqk8BkD7/mOGCw375xdMAtbqIqQxVURfjqeRChOeQozuIknMgJAo4WgwEeP5Qd0IRA3xz4KdIM
NHTHzCNEN09ozhqXmNHFPjsU5AZMgKc2X+AEDrf1kCmzNfHkGyfrqi55soX5T2kuzi1NGHaGvI2e
wuRwe4Z1uZ10L1zmvbX1+5X4w0DklrGxrhNVdAqngRvGd5R7hNt51Hk+1LTD6wooN2m7n/aXi2dr
pR0U4y/tH+niMrnDuvpuu0MXY+lATbLrJTDbBcv+33AqWOaQy/r6oT3D/cp+zpotmHSIj44v1+1w
5hfn+TzXnYaSRLiKxGFAXlKdCefC98LRewl9jkIRSHS0bNqFnY7qju7lJPCqXMLZwgdT8PNj1GWz
t/8S9+aiygP8Ldv+12/gOKDHawNZCXbBF7iw5+SsLBvilXbBqkcVviU2q5dP/mR/Ccy9cHXmeCgT
xiVgL3FDlvhMO6dgMEu+IuOFIv9B5E75hlZDLpZR5cvo00zn4w+0imFdoYcXoNO6l4afTsPRoOXv
MIfHR+y2UjFuIt+KBl2wxmCxbss7qwgmsXvz7Ng65OdPrYj3yrzKpo4RbE3dXqAhYfWZQl8sAQt4
hN78bhgPjyvgaP0dD1CbkfDhuB21TXdRWnvo993QL8bMspAoo68APcatC6mAbFC1VQUL6Dvh6iRz
esMJVFKrojrRLzwd2ysS4z8U2lrHB0CNUMoCPL6bIXPlHMTT8UwL9rK85e8JhmkOrWHpvTwJqFwc
N0hjUBjySFHaAd9splEIFzUGr7W5y1hHAoDdqHoZdlTU9vyX7WUUsadzULeYy30GA/wXxMn/p8pL
x+SDLY8USweTOJBmZZUKPxfGSzXH7Dq/LW+WPWRwRWVQWACz1Yo9MY8iDoAEej2H/StgSvUhTLRy
5ZiPJCnS3f1Vy3DS7wx66HqcEelMokZOSModUNnsU2gPEGeeZ94nq47j8iMS6HnBCYqK5YAvwhDg
ZWRP2v7gNFQsTFNDVNemJcYO6lIk56eqFqZ+vRr6xmS2SZuSN50EUKhcpKwrp0WLmLKICgTDoneW
Vo3g1BQZlPOdZ4QEO0aXlinw7mN1Y7JXkweQGYFvkkBdXECzCzlphqrwLC7cE+xMQJDrljH+BOqO
6rD3gey4W58L0BZ+bbNoNUpeokoldQvUrlvYXVaGnVqkw1AQhDXhF7JZYNPrQXt/7eCw0LuQEIN9
k8BsURdJhNPtXrIFbxFUIcxFLCzjqAPcLbUc6qSJIy3QsxGz9zMkp8bnsbAGBqPB0WnzU+45N/th
DSOx/lskS3j5PyDdnxRob2lgC4uw4qFd+wJu0feP6RY40ymIHUltrW9eh4Dwcc+OH5OhxOcgc0/k
QQvmkMTVtvGlUZGE0QoSTExN5W1tBPSMVOuhD0iD9SPKnacElU0liA/idQ/sRjUS1zeqV5AV0ao3
QoKl2PAmzVTw3uWnB1d6cOoSzX7uxRIkPow0SOwOleb73C9rWhN3SgFfED8Cqx+f/Vvdf8Bz987+
5vM9q97/bbT2Bi24xLefR71gDzNO9WGDeriIP2wZO+Mg9tnZqoRu1RMmheXWnLjmD22jinI6tqyG
bM7udjBPJ7OC+D4gCCMOftzKWzQ7ohx34CFqMSOD3Fch6pujSVpepIcz6/P0rNfveF7Mx5g0gI96
HBfHtYuSAMDhccXx/Ic/vV16Eh7r73b1DeJM/qYVtd33XPMkVEFHk71Dqr/PFnCC3pYCsSFs0NYD
bZEQHujF7Zs3u5pSlttI9f/0CLup9UhfedKAViWhbgumrhng3m2pdLUBs0hLdFmJc54dqWMCV2Dj
IhWToPK2cf/v16k1JEXiqL6W6w913Pny+DECfRahSOZhJirXR9enbMS5ii4vNGcHcd3FddZKbxnP
J0KIVBpXTVwZDdeh50KS7O2qm2O1VxlSQ8Dk0tc0zJSJ84OXd0Irwv9hrpdvQXXUaLu4Uds2wmOn
hdxZXIwGz1E5sGCq6Ma5H8z7AN7FaG2gQ1CuCDhhjBiIzHSIQ4rGbnVfoRcAVxvALR6EnWN+iAfC
gMN8ZnKuhQWSmDzboEOQcBhKnxv/i81MGWWm6ETmH4wrJhcu1PTA1EPPavrkcFs2hYKITmwoUYYS
PEao7jnX1SQJm/mB78yzmUYWGp630f4eEiDHmp9GDPOciYK+zkUqtagzy4dTKEICsyOwlQUOTtgf
W+3/MiE+WALTByoCkPbRKL5FBKlFc14mg/R+e1WvMt/2A7zJN9Wn2u/DSztbQtP23m4L6cloTmvF
tSozAncibOcEjUNDvZloUVd0hTkRWUjiwXJiE3R9V8fB9D97KL91BT7wY+IfMWV7WXxZID3zK6c5
KcRZfeKY+TteQAmJizB0uf62a5rp9JoAXiiHE8VcqjnWn9JKfeDmdW8WFh6Ga+ogrM3iqc9HSuKz
a/t1/TcSIMHEUVchqCH8iTFozoXsdXTBZJ4hJ1BrGxbGjLRlnUcam3A3yUjMDtIiDBfDkJcPsHVF
Idl18u4p3MxF5SUGeGcvgx54hGsZ+Wtk5b+OSkBoSzmDifspc/01Azz0rDPbNt8gsJFOxHTH93gq
AxlFGpiPsLEOcXzsDnubwOMJVqNWJGuO15wOGTsqL3nGG6Q9Ya7pywFgEG1JvZ/h4zp5RGnVadgg
vjEWNk2ecZoROD1eiD9AV1UgWvK5HT3TiS6QPdkKjchLI7CpSJneP0YDGwColi/CNIKyHCPiDPf7
7hYYvVvs18Jn2nYxSqk0kNuyhZJFh3aaHlqvBuBZuwmtBjWzfQwIPhhXDEC67tmlYaL4sI3QVTwY
YYQBAo0KBhcSRrciZ3b9W9jRVHdLLGURQ+bNOwsw+YcYos9F7CaB2m2y+i3LsV5yyS8YFM+NOTwB
Sbn4yRwH6tVcYtMsAPVuvEcWTyVqMel/xyG3nALJlWJ5hc0+D75VcYhAIq1G2rshm8g3YC3kQwfP
888Q8gjcIC9CjBw876nRrE4CBIyvYndWp4VhcoKtsYfF1k+GfxgDXPGptOTJP3QDSGUKyEVBiKHk
TPojrf12R16IqVBpJ3cpvWF4tD9d9C2ahKmBP7QnbuZ7r4gct1u8fJffuCvWQHqV7t3WbWq9lhCs
soFeCpZn5CSpqDE/LYgdasxnuurtikPK0w1UEQC2km/krhbIRb8J3Jzv/9BWgjs49tJB/H/uzMUV
Cvik+gSjJ03uU7z/EKWsLlyRsfX+eqcU09wy7mo8GUrWuuhkt3bs6YmnAKiHBh2Lt1ptzkU6jGvX
7NmKT7etrtHSRhqdvIa8gU0G6NiK8AhYWTHP9mIig7fddLiX8gnQh/V4Zqci8hvtiRz1Ep+y36+b
1uvbKBKQ7LalX8YP44fF8Vh9X9mAtFYPA5yWSW04Cbx2b1fUXcK7L16iBrdU6v8EYUAdGgkCkoHp
cKBlqgadGnQAnBzql2EoDH8KTxIlc91fZY+TIUPvlCdAABd+1m4FOTr9kLN8n2bNapNl/7uDSmY+
zHP/UlCZtTTH6epW6d+TBgd/7xmilJM6EctM99N1veE9DUbZO/OZ5rQ3xTK8eOq0MO4fS54vHWJi
NeqB+M2qfWxZ3E+Y0bL1BEXSDysf5JKtOhuXGV8L+ZneOGRk32WdHhOHG0nr+1Gz7+YoZgq+L1Kt
V02yThuYekKLVAqYS//6Gr6j1fPWhKEN3DFDUph0HHMg3nu/Vd+UFvmvo0XX+GDNCfUBz7nJYi+G
fzp9BkO6Fz0+QAUxkhRw+7gUtOXpiStecqctWCew/9DHj4wcqhZtlyrVGLgK1eYQ0zmgiDx2K+NG
2w8uXgJFiw8KDd2YR3JV6X11DXMcVXqNXhIf+nbczcOoMWgmAJ87oKSBtYV+FO7w1gHFdTgPrF8F
07ml0VgW3nvXhWwISJN/T0TbyG1UV+X2e7LYeGokqNNjor8bp31Enk2XJpwYZ230lYvXkkztPJkw
UuA3u+kZVSA95oBHnZCXJeLweONHhnbw4uWgFVGm9VV3UxzEhbYTPu8GaWvJTbW8fNKrZX42xTeb
P0MG4CiHUE6U3kOuZjdf4JGdC6ejK805lH9ebxMAz9RnEfn8Begn6Ak1ivGKtXMU7OV6jL5lVV56
tu9FRvNBHeC4rC8lh+vP//O7usTceNtFLLEXcNYARwX+eA58VNrbt1di4v/9UdkRHnkNmARdYcCd
w4KxFZAUIDW1MYcyASb1B4oc0nt+Uq6hV8O1HHiTjl23/GaMkGL0U9nHnHvSnxqH+49IvjIDpanQ
zVJpQKApsihF9bMXTTtCrwbVrwEtlYaRQj1wW4kIBVy48v5VQKXO9PRapt/PdCAN0iuPCCGsuV/3
DHPWemhTeoE2vMqmlUDtM/TOnW2DzouS4w5tR+rMdRMwYHQw75n2MFw8zFk9mxCpdFLb9LXhdJmg
tUzwNeYwTPCKmIfMv2UuhNHt2r1j5q3qgedEVz0W2D1v2EWCNOaDNSIz9SWtXNhYKJmrtDwsXjlU
VWFZAIttzT7z/2QrN5KvOiFp51ZrO1Rt552Y1E3HNfQ2OHSs9QGPV6ArEdIr0cMCgYx/tSHKNEtZ
21cIXOa9c/EVeumOHXTATdqnWlvVVaybugdWrrjWtfRDX6/Omau36K8YS5b+32OpATzo9LuMzmyL
dIiIbOjFEPFNqqslyxSNjF0QSXimxZjGaZo/ZvTQSfUJsRpqpkicsdGaSZL0DKX9lH4znfbZ47Mv
fe8nuOK5EPLQMyAHOAqCgmBL00aeKUeyjPvee7g1eLQdm6zXpa1E8FNAwdi6+ujcZErMP+yZylxb
P4D0wI6oxKM0mpUtkPDDfSIWYdJn9u3KQUkExWFPVeS8ShHgKSCE6uEkeajEJUhOUTPrBvX3UAcF
2RF0cQpn3mqG+Vqq0oaOw7pQ+uhilAX7n0sH8oxqkZAf+cpw5U6pK8xVl/X/9Dl3ovgH3SUEEkAN
aqeFDgPQrflLMel8wxr+H8vQMKGbtaI80z3s4vuCLG5iKc3vqenKO0HcgTYQSv2Cyso1O4x+oxg4
lklwZFlsTAsDYiUgewzC1bWZZmdyINOPUmoXA7OFUwe8QJUf7V8dPOhiLEi1TgW7vVpMIlooRpan
ImjyEh8fu2fOh/JEkILLORWegvzynqmLXFZ0LvRhQVxmaugEhZyBJbRHO8JgE7TycUTFt4Szv/ew
/Qk9+L6KtiwO6AmzNB1ZFmgOprVBod3aNsYPpJkvuQFqsLYoV6GwOP7YkBZ0wkS5YHeVZX7Bu9IW
xKvndVqsov/Vayc7TVpUSfnubn8gKp5M4whdtxqrxSPFSAyt8rf8s7e51ZDMVfm0YQRAhVQ8LTc6
9a5lGyf+u92SgSBPVDUF33DRVHvDndIkp75h4yynqByC3xjieHkRQxn/qF9YNDSKHM9avcoxoUCu
EVpElFHvVk9W2U3Ryro5WZ0PhctYLqZgwiaERQUQV+JKrmLdbtr/KbTZ6kUXUtjMqA2UqaZ/yU/Z
77+MX+lSCW2rtMq1zVntRJt27orG2yMZaZUEKzlUwSZe5Gex8yMfyrldsPSZ96LcPvJ63/MrIIGc
vDp7IDJYrdKWX8FuvL278vDT7aADb2jrjW4baMs6ZhsHoB7FDbIILTMrBxyKN8Io1mSYw2GrjREc
mv7GtqElXmwZLR6yClpkeyWmCDQZ5S68Lf+gdKT58B1w3F+Hx4KDKYWQ1t4oUYR/qH5w4U/DGjkB
lo/iDUa+bsT+dw9GN5zVDoJiqyNbbTt7e+gUvJke4RpDdqmTk34t+HeNb7iwoYPc79JYueGturto
gGT9uucMywMvySRVV2OvHgMUZ+EzcTQgdfkuKsVEWrmTKVUsKCADALq5nHlOuuzbJXeYN6XhBRKY
unujBui+NZv4IEwDL9HtYnOD7Gyv38L5YimKA5k4DLvacSTAIsp2MDD4c7d62oliAXcXCPgPiyMv
UpucJe1vr4/7F35HAAs8asYYttR5AteXQOiwmL4W41uu0PlWQgYAYYMYEhJMfoIKj8TWgCPlgOOD
qZtdLE0BX1VAVDuT4U7ZVzvtI4Z7l1elDTjKKN4v7wNTUaaPyPS02eMONhV7SEpD5E4XD8SlfpQA
igZp9xmCao2/TMKL+67rBQuq+RY3NGBpbiA3GS9sIoqY5DzrXVgrbOGcBbLP+RRCaGobLbs4hVPt
4cnZKYNLXmvOW3Q+sSAMF+b8w5gxJZmmKuDkrIWXCULd3rwIrwMKZlLrQGA9M68IC0ryWZw+Gn/Z
UiSbSudGFEy4gzV3tpQClA3ttHpliWxDFS9+/7Ie0y+m9QhTztoyQY+KgmF7Gg2A+9pVtqCMNry1
+IgGFw/WYNKhymFp01JcjjtVePhThNfReIrjpcY3uhrAKcoHjL0vK8Vk6LKhh11uGeLOH759VRHZ
YwsMW6iY0qSJo8BIHwXBSXsD2b/uySItNnthC8u1H5vRkJGeHIM5/h7SKmPCXFYhnQpLWaX+4MgZ
OBjfeUknTTUixjcfDWm4vcwhWcS6oyVw6syzHuZgqi7MlJ4nGnNtCSssnsZiSC798WZEDIBo3x89
IEvkZt3V/VkrCIzEUp6ZhBwXkgDEQHfm2oe3Kr+0xIYg0qP7Ni4I43Z02GNDwHVKCUHPoc1of9PK
SLgeU9uK/c5gy/9HBj/3pP1HASZ6zJB6uO550dwWYaC0qG/rbaSRlIM2wfJvFvRT8ujy6OeOIVtd
12VAhZG6bmnu+ZyZTq2FCRHbJ1kE/raR1EXMtwzyOM8BuTHgBSSsTUebVxm7d6Eevszp663eZDKZ
wBq80lQjuV6qTBuz1eo3K1L+zHHC42pha9c8cNFQXJE9iVl0Oxenpcp3zRA+y5SCxE6hBt55o+dL
M4jKGHoT09Y0wxTYHF+p3BfCuhi7lUet9JMSXhQedqWvpnKNHiPfqBsIrM3KLZqwvLOMWWaNtr5X
FdEaheS/ItgnCJjMeQdYkbusB918imsbp9VddXsnB2PgPc+Mf1wuhSCUwh9a1lrCQXgiNKxKYJuz
TCpBxbTUdayX+mlximC5sbuxXY2Yo89q4uAb4S8dwXkX3hF0GBvBmKVrBw+eU/4xkF5C/UnAzZTN
PimM3+fUHA2Ff0OL5MYFaACc96Rc0Q633yPHUyx/KEI4BfGTEr2I3RLXrH9P35wWheQ1/CYauNIX
E7M3OEwG9TZVYfWtWTX6jgeKnR2R0gldZ7BP+tzDcNLZFHtzQF3jHeFRme/Rews1oe4QAWJqmLPa
l38gNfiFZa8AA4nEAl6BPPKwb3PbFVDwjYm9cKh28sF+09WRRgJL25XbB+O32Ffq4Iv708Ts+QiR
yDgQ6cZKQuE5GfajUpRygA1UNz/FVdoyol6IeOVXNd+c7JMXFGwHft1ugUKB0VmsJNY+6HCw+BrF
dlI9IQFLQ5+QDRJdU+lqf9Zva9OOY1yPmLEkCeTRHSgEMWul3bnMKbdz4y55aKNM4D9xxrPNgCFX
E+Ex8M5XknMRLdwVF82UAYOn7/Rw/yzefc9Xh7FPN4uHhgas73hYDgkGkv94V+gxKYWBcH/p2IPl
XzbY97R13IWKWIZ/9sp407GYQeyDbeVHze7CP0lWK5uckm2lx+eimKv0p5G2f8mIfMxMF5H7SAzX
8LD4FwMkikxJYqk0bZa7noXxi8hJVWIcudDhVC6EN+EeyIxUI1bYtbwTWzCYp5TTUHPy3uVwXUj6
aMCc9rDlLUDkmRBkbQGH43qHFHMoh+pdiBEphS22bRrLAQFGDt4yOuY/0obroGIe/UHGHKdmzW9A
UwQW4BXgZWVPzF9+3WaVmoU4/PHBv6CfPN3gAbW5kgtfxPEgUPY1sNQDv4LCGl8kAya5XTcmZSkF
KIzNCff3XejrAye7gCJEb1wfXR6K5GoEJgYLBENViCXZIwhYNfMb+wWbg4sNOhR3u+8hai169++V
Zdd2YrvTmNmGQxPplxOnltq+4jfDm7LYILK1qC8a+HJaTcRy8Vp0nJIXnVlvKqFoDPCx3zHOGMHS
QayDTIqlhANWL3C1ojaoE5xRY8NJSfHXCtXj8qGZ3FvIiB4vlXMglkl95e4OUQZKs84EyVbuXTcl
0yJOXPfuuKZOcLrzoB4tyep01Y2+rfTceWzx60GgK7bx7FkgQ0WwftQhzYMwlUo+rQ3X6P4dsdpF
bHeFgFnEJXogDUMK8u8ulDLHVNxhyIzVihJ+iShdAME0dTKlwGyDlX69agpQOfVxlVf8Yn3pK/Om
CZRLEMgM/hXFhcF3P/74nurZa4XGanG5SRMvU0Rda47IufTIopBOaJlst7LUcu6KDUa4tuaxyclv
aj9xMmrzEtzzS4VBAdRX0kAzuZAtr8/KQReqQW81B47H1fv+qcDDS59H9ICPizJ2tt0gOR2EC3Jh
InV/NZizRLnA+ekYk8MwvldEDm/6WSQTEy74V+ZPmBoPRrrExfNzO6HxVZzBiWri3/kkAk85PjSi
PtqO2lP/ZVSzRxY5cX+0r+HRGhTGHZD7cRxmXbLXba1VfZTMpivXYPryR/wROEGvlqOjns67mEJj
YObrHxvOU/ske/J7ruhPtuZ4gmt292Ysfdh+3qL7owzcVOL7ZBcdwdXMDF01fOIAmjYKlbyY9X3P
Ux7kBdc54CxioRWR67jixQPam18zdK77yBKPtdaaz2rrQofGoSRcmSMCtPh9JcQg0D6bB8eBFvDU
ijjL6NfGOlSsMSC6kg6I1WeKX/GMqQbpcl6hukUsWh8CRWeVaPcniV+aai3xj/9MHp4OdIu6JyaU
KJWPi0Uh1DVCW7xBTalbC+XnHxrB+2KBbVEPFxusC/bsvzmhBNFdRFvuJvZyoQBlAWHVBOHE7Odc
lC+9LKw4YonHYfzPe8OT2Xigeqd9LOSNHyNM+eFixSbh7Jx9Ed+3i5ZNo8qIkOOE+GgLnozE/wMc
WiUFv3A639BwAuVCT9ujFzENCr6Wtp96knHPHEnr99hEv2CAf8z+cQ3Lo2I66RGWgfkdNyC2bulr
a4K9Zk+2nVbe8LQwFtIAAqR9g0ZtjyIYI0LAjkncMWLWBs9opVQW/8VGS1Gooavr+b6EZEr8lJCE
fuo1Op8qwB30WXET/JOxLoP/BNZILjf2yk9zW6VV1fLBA8UztVB+lTO4VFgnrzU5Y2mCaRBL+4gD
IPSTpAUBVEj3VM7/zCYAXXw9Mmh5DrNlXr/L9jb8JXr4vbmmEi0AxNxd4+XUglOEeg8KGom51dBD
d/1dmoeASbWxGTJfWUgKwHzD0hxB4DgR7zLlDPEXPGWGEgyIq66L7Imi1DmU6DR/3GM4iLYGAoVI
Uzu/35wWFy9B0cXwMCnHBeF81E+eVRm5pnIffPBLmqEAI30eqA+YfHjxt2UtESql55lidZKgrpj4
EVlyfG+ZjAvGSUFNyhc00GS70LF7pwee7GdieoSt+A/JVvQEMdJlIfPq3sjkaxWAcsW1bpQQ1iP6
jRqMgxSasgs53o9Rwn8OJMQx2Thvw5SeNAfb68XcAwTLHokUXL3cmRkY31vUob33JKjQi4sN6oRi
fXOt/YXrhRYbflp36RBkqY/UjpoNwMiLDp1X/1Nw0KtrM8gnL9EH0IcpDolCwZXerKBSm+dJ4L1x
LyWfA0B546NhVBZgeI4cTCpLE54yTo/h6dyc5QOULTfb2ZTsnsYBKEwjjacMo0UE7RrCgNFMPLlN
4W9i/ixL6zDAVRIV+CL8Y7b1cuHPX3N+YIY0GqD4KbTo70DHBR/EiKOtX3fLTwLjhC7o8EcfMB3j
EeO8E+7jrxkLj1SnGGXqxHYdDmeifq28WeKIRDp4F7n77m2diDiHktv+iOi7TjDeOeF2ceAV/TVZ
S+VLdhdgEf3xpQNyfDwXHMe0HjIOx86+KfZTxjGnkzGv6HSJgu6JKpvHwics+tced91s8oNh2ESI
RaWK3ymcNij83x+dxe7cgIhli0YBs8GFCeu/1PqrLLER1ozZmNXA9P7tVWKpuo1TWISU50WtTO1s
/2OTopmCZoSGON6nhJW4TlIqnl6Vj5OIlF41gdofvcv185qkrIjnhPNq2cl/GtGm94NY/dt/aBpX
NrGij8Mz2BSJ8xxJbEnpidm/Bqkzp0Ovf3hjkjBnEQAgiZJWtIQTuI9OOv96DglMya9kOk0NpVjE
6T9kJxF6vNrKwzIQO4xImhPbhzwZljIwedGIYxF/VrMLFCCnsNwoOYAklvj3IsIWhHli5mwvuSer
dytLz0LnEDqIfRiiAVKgUO2nq6P/Nu4lrtqJhNnMJeL+tBSckxM2x/X3oPcicqAiBmQE34Egss6t
WjX/sojRTmsoOHKNLo2KVUeotQXSAh2lIo68SBsc28/ZLsbPxTLnfGrR+yrvDe2p8E+3NdE250hT
PMXXP2N5c8w+85Be3n2uoCcgjaUzEyBwenPpYNqKblGADu9/U412C8ckIJeIQ6rPhVzPioAeL/cm
a4KawODYZEosz3l6E8zUZEbn7rYn6C2IGiQyYHFjaeEiYLEbXUrD91cORT5YXNScwiej2VGtVTo+
K3d2u6jKTcxTxuWkiwVSTOct35i+GtF/ZgSAZ4MdCep6mAHmNsPaAqaV2+s13Z2RrkeJnay9M9tx
lba+r3EsuSXd4ajvvxMkkuHrjt52qMINr42mW8gHFAzx14CGcAtUID2NFslca7UKwhSl8h2lpWD7
sJIGNoju9JZXUagKz3BnYstVbL50DuyHjOs8tSGSW6dzmOOK+nneNm0oiRpZ6SaOmp4l7PowSQ3h
rGsN1x2noDoksM9prtuEkwr4ziAPm8bUH3BEUkf30aoXqEHZPiEAN+G46iV8A+HRZDzbE77lcrqE
qHKY8q9bYGBziNeORFxrFdvT595zs+dfzi+aWYo2bLPXGD0sLXRhza/7qpIY9pf51xjbHhqy0fyQ
VOsNwnYUMCRWcoSMRzCYYAKvyj9cZzeoAVmEclscV4sVg6UTQ2CMYByZwGxjVOrWkc9Hht2rQp3v
+p+LN0PRDByDnnX0UVVw81Bu64IqzRXMhAiBy5ykoHbyy15vm7AGDL1Cz490FRhZfUGERByDq7gt
xyMpqb2SUpubxh0W3t6WmNxmkEPj2eUx98LLahxYF8N5XGpThXvVQRO9HakJpVkdE96p/6H/ka8S
jGdswbGVlWAeTSWGwUKFyw/rnlA6vT5xXvm8mf2ltU1E8uIWKJbjJbw/yn6GQZVusEqK2AgX4phM
avjt2gr9c1bi2BLNldfXQyyb7m9uOtJxCIRiYNN4pP/KyeyFsV87sevyS6pFnzhu9FL1YBENLUPC
SiLPAckykS1CvhWMiooggiDSsWe9AXDABEkjtATp9W5cU7nlkalt5AHjeg+nTtSy90TQ5AJI/RUy
1U0YDO1AhSteLDVoLxh6xQNKrCachuyM7PJaR/iCk8xyx2i5iDv3Joy8JA+/zz5VOCznFeFZFrPM
wrxjBT0m8C9kA2cJixnWdtd87Ks3K5BI4rJ0CI6VGdwpp2S36nPd0kUt+FPYsSI267MCt0sPcTLk
5k/R6AdYsrI2/nBBh5P1WbvG2qgWe4ftCiE57VwuXnv7FnQ21ZhjJOZ10ox2e1hmUBTdhch6IXXl
U77u0gAVXiGLsw+b5AC8F7ouLlM7iqC/vHtSX3Dg1EtQrtBo941TH1L8x+++o2e+O5VMJ5U8LBZJ
nVDg50zBSe/lIhUH5TaGueHiGdmSTXeKH5tnX2Z4grKIxCOG8qZWYXtoRTc7FCB38h13HLl7dxD9
n0ptKXGRYWLZlVZxTzRi/ihh3P4Zr8T5cvmo9XEaWi1P5xnghdkAtBY7wpzx07ExgfSL1jOGQzXm
M/w+f6C1pQ2j9HKyDm3VkuU8lH3qKljIZrFM90gGwPsjNmsxI0c5J+U/9mL8zhbSQgkBdNj+aiAN
SHwA/ba4YXiqtNWOJ1jEj6KPd7YmggxxLuf1FpHscg4E5eX1nhLFNV5m0OFSYQNDfLEMLR7Kz0UY
3TB7oJWH4iPZ8FjC2qiHFLUHJUZx+M4wZo8ZtEOSQ3onakWbeCOZfHl8h5PsvNjDhWg52VR711/V
6x8chgV1TGDRp9MB2wr69tQmADcRI2Uymq4D+h7ttMqKDZ7bJzD3I55Uu4KipBRxhucJIV34MxMM
aBatP/rDdhyK9Rkxog9NYBIu7G22rQm/S6Uitu6d5fjYV4XB/0PBH5o/h6g41iD7+GDugQ0wtVFS
3Inp//Vn6LoLk+en0FOb6fAMrSHWBo45CfOpMSPMV7BtPfkxV5Ttp5RhyzDGVHCh/d8hnPIrpyBR
4xVjxNhEq2MgVxdk/ehqvYOM0FxqFu2d7XigT9GQ6JKj87+S7q5Y8gj8qWAXDnawulwfRT6q/OpK
XRqAaAlOlbpK4JjfLPn4PRruOLi2gFe3oQWpkKINZNe81hlQiNHmKbq+D8xwkzkfXx3aS3UJAZ5d
bHIPWvV4ERH25Eo+FQRDd9Rfs4j9VorsTLEQjL5YNi/mABlWn6PKQrukjWyJBd3pEGA5LvN7NDpZ
auTrLk/D+DncjzHuh+lq6bUMrWHpzxdlSolT3KLxb9BeMgj3qtff84DZSKN7cl9zeya2Wl05sK2S
e91k+Mg1uYF3OtkG+qO5cnnK8y668H7lx/Beos7Qw5IEicibdWOoK2OW+4j8+sVQFvhY8mt2USqO
OcsFBCNp9MnEWqT/p1uK+kFhi5XtdoOxGVZ/9CZNVpL4MsV2ec13CfquFmjfWLMuHvk39iMM27fW
GCg/57Be2TAh4R2cpgVm4pyv73MNCzaxySRbX0VN6PXzykBmne4us6+KaTxck9xuGyr+tS+atEN1
bBgNAJSGSSK3MnL81n11v/AXCJlhAYCLLQOcm3LVIvOS9nKFDdGQZhmMGePMnX/p1/kyZs2pmXc6
fA/hV0HMMDVOIIxVL8FFkS6+XMSeM3PiM8bsXwKYOi1G8KnttMqzx/UDrrIndhFGW3IGdVdT0o0O
e7GyikMyp5LUOFyqSkefBKtT2D6VFiYR8xe36as0w5AmZDzbFi1Llf92mHUcDaPEeOZsX6M0Efwm
ntqb8ozfpJ23Y06fT0Fv3X742JiYMxNaRHozrkZfupzgDSTXksKV3rgMtxRlXvUPOB4jdiDB1Zym
axxH6dfcBU6L8mBSgC78pw6jJ11UxGdRt+6fLbpU7n2NXl9wPhUzK/jOe8dNz2biv+0t85c6qYRE
SpaUn4OnKh4GTr2PZFxD0o+cTKwDN8TPvr5XQkp7TTc2Kq6bVzoF6JU1+b5iy+DvBfiNs2GWCA7f
pS5bDwyhrLKRQN6xD0oXzTfkmnlgxDVtodbq9b/WE2gXTnS9AuGd2sBq29EPD0Ou1tSpONwCva6Y
oqRR0DvO6s80CHWTTbiXVHcwfyzxT+gen2GZUHDwokWKJpTEYh3YxB9FghTbPVy89w82KYRBuk44
6ZIjEfFcX4hAZsT0jkIg+0EWOknkylDSzKkrSC+QufAJ6rxIZcXRjNyQnQcN0zT06UXimtZVhqX4
btXEdFsmImRW90tOsFCORyr04edbqDMGQqYIuasljilZ+QjB+nufoGHMXGVSluCk317eiuJSlLsh
V5WPM/TxcMsGmkOTFsaFk7/+OJZPyuvs01zcl32puPBygxyj7P6on8fLQ1/0rnBCm5kwrMjkEqTJ
oMxuvqqIMJ7tU43I9Lcm/vUTd5fURC7xaMPI6Q1tCfBQobxBMo/lUN39qXwE22wqGRIYkEemA4zd
OfeFxglWyOgElxJs2ADK3fgfTMcoP9dVyxjw7kV057rPx9zR1UHh3K8pWLEeRA9uP/Yj/KtavJhI
1YlcRuXcjms94rfZniVi/5I0i4rKRiye74sahnOEaONRnx0K/DpxGM0RdnjJ8i/+6jAJ6r9bkqEi
OzGEwsNN+kO5HITWL33BYFyssz9Tu9xpoLAuxSVkR/a6u2kWQlD9/LSJ8yXaUV7rmFC3eRhcTIjT
3m8tw/w38trWnVEH254Ql0z2xO9zVhm6a6wS2OrICXZOaC+dgH0I0ekPftanq+RLDjl89vcQ7Iie
B4TTmymZ8JbudnosPDDZ9tX/+Bvp9HywZmecDRlzZ283foSVRrtAbXQCzwRCjgYz6ffuZZKCHt5Z
vU2ywseuXHWkdFmFYyw+AdkRa+dcK2W28BLGhewg6C70yWnU0aIQHj+PmBqWdXMUVq7Wypa0iI8Q
vU6psJwiwHFO4cKBGgNuvIBIelOVkQmMqE40J8eZ8fozvZxhTPVmlAITEsBeonC6KF5KNEz9E0G9
vXhSmnNAZNtWstIwy/4XKMRc4mVzraL/FTuBCaC2yy30meKVD91caKk4NgqP/MpM8vmknZbtVrBH
c6v65834MMJ1+zQHUqIOzf7zKTCB3i4dciIllH5qUx5YG/Lr1gJdz1LjdWSKwn1i3DJOahQ/mD3o
PEfk7fU1+ZB9f5MaaDiSkIirT+jOJ1WHL8m7LayPPq75Ob7gUNVtwpMavXfW7n4s1+1gzBlu3veY
9mBTXFyczf98YDlcrHPJGSThWIMumSk/WyEuB3wABc8PF/a28rUbXuGZALTuNCbfd8650gwqEvu/
a9tF87PEHngc2gUUIF9yuSiQJNwJFHgEh7+jMAnrfaM3vnxSZ3OY8Cqq8LQBMvddSKLgx8qRnIP2
ggP1jmVobaXiVHfkCES89cZfUprEmC7cR3wuHIOpg1LMgiQmnvUPNRleYqoQ3T9jvpQV9t8l94uK
8r4qLh4hsdUwaJPfQXZ8zRm5HYz18Q0ZDHgbDjM3eU94Zr7GoD9sVPlI9h6kLrTYsL7fawmyqdtx
aDZOCHPqkJ847W2MVIiLTDncmdOUjAIGFcY5UI+BfSLm5VcSzNMCFWltG2RzDK7rZ0FI/qg4peig
nyxVYkBF7BTv+n7wW8aiB3G1dGfmb6bqiu1kkC0jTmuOOhkdaryITxvklr6qYnFW1xjdMkkB800m
F/k5Oll7GfEQS2DzxlbFsXV1tXMAp3iPlTBs5K84FE2+K332qyEnNnxNjMVTS9Is43vHCPF52nmM
Q7vsb6g9IVKJD97ofQ2Zptqut8v3IvXN/UZ4ia/SfeepHbs84+r9siVKQ9x3uPKAdXoAxovRnHOZ
3bu3y7PUDWMZ9XCf4diQGFuJTMDI+TejT31KOdtOa2rppiaM0rNKv/Iod8MoX+gwHYxgbASf6PHO
nZhDzZsfc5/W3l4j0GziO1yOeVyvnwePxggZi0fIkBdvEk+4a/0+3gsf6fypBkncLHMqYbor75mM
vusiaF+qKfF4IZCboX9Ksmdt2OOyhcqU+ioL1y8MMSdlTKYAoXB8E7JyeSrFiZl/4O2Xc5lDLz36
o+LOkN40BnBN7GneJ9OyoRIGdIg8+rMoqDYOPpNPgi3lP1/ffmaZ75e8uy5r2olYQIRot3EdZ/XX
GGvwK1NA7wZTqNu9wrQ3mitaPip+Xay38Drq/Q90WO2JG+dPm/CLtTULed0qRGhGsbASDqSGIgiu
RK9BP0PUVnozclVknhBC1FKLssBOeIPAk5ZyUTMBUK7DWAZKpOgQNrgQhlRACUnq9fjtn2v2rFFS
9ZvodxhztHIrvstwaiMdLv4nvYybJ/aMs6gD/SmZo6eOCBU+eueO6eIc6akH3Yz/BTQgqoLO4T0Y
wHZJKNkbGWKL8T2lTXkEHSjpJh4d2k4j+rNDQqEmntl0Ha+ihNrooe9eJPJGMz+vJZNEMpG+ueCC
O1DKdoUxwYVa9J9Raa2+LhD1RxG05N22Cx3VhyLol6nlaNgOgADFLjz0GtwUFLdeYuv/n+ws1pZv
SWCN3D/dqG2zFVjyetzIgRp4w7RuMWeuBl2J/KKOdDPG1R3Xg41XY6JOYdbUqpGdFMledU3Xrr6r
7CBf2hVtt6cynhLVSeb3FXf75tG/MWClQ7IJROQ+jAWR/sV1BoRdRQ1+PtYUhMRemu4CXQyvkYCz
DxMDzxb4nkxg9XoVzh776JDr3xR+VZdERkYNy35acUvKODCGieFV2wXRZK0cu6wo5QvqT3NAmEAm
eqvSGhMEwQUMclJ9KD1q58cmiYVMOKp7WZBDSb7MIayhOAKMioqkH+84lUULbbMRrlFXbIiTZO0W
aQH7Rng4Cb55Qoxhhs/q2KNTEKAgW2W7r4Li+mFxt1kRua2/vDIOH9dokG8wYqAqnT5FQ/Xyx4j5
AyWtEdCZQGxbGVdYOhlh0LookOL9pGauntlbtvPDHRd5LFiNKeSGw/q7xChikf5pPCnVYGDSVe8/
BKYs44zZ2P9qK4XUxDQoqfjK9LvWy9lQmuw94W/xbnhgljtGG3ZqGE4R6HKdpymbl7c/UOy1CcGO
yfTYMWewcpX6YaC/GPgTBEC3LsJBVYdPr5bg7zqlbsuXInWVxgcAVVV8GkbpRWDTzNnznFsGLMiO
83BXkiJz6Ccv4aFpG+0RVPWhIzqQuBEfu5Np0gH4JCQuGvySWl/rVWxSrPQEVyF8zchViazn5vCO
RyefyOdwWNEijysDTzK+iiN0yimXJUolCPIeD+6DBqMSHk4DGZ7mO6/40x64pHN8D98vpLOBU9xx
QpqqOXIzeeH5Yk379Ij/SK5M0RUSgCOtahiW/thuCZuP3hz2zMWWGcEiWDCos1dAenUeIGF+33q8
95ZQURwiVDEokMOP9gAQahEQA/NZ9E53tzTWcbXRYMuHiQLXPx1B9tQAtSAxipAUkuRlr5hR0wsK
XI7JnThi6yQC6QII4DIgL21CCdDze5ag41TpMVPzVi9kPlBPSe/b0yJvGYv9qeNmQTCxK0jr0Nbp
7cokTbDj/aJ1J5VCaotg3i+ZBGruW/W+quSQ4eilByn5t24zdDhIfoBa9H7CoWreyNakLZjeUW/F
1eRZhmvvOHa9MMyxY1SFmDPLw4/YMK36nqpbo4FLcrOFtsxftUfYACrYC+WHizSTnGZ+lfIf2wu4
JTP754jUMix9TUOQvzIJUJjuNxE6CUKsEerPwp0Xne9cADURTmLaJ4mSnxUir5JK6KIQkqTU63fJ
BDF0GW9Fez/xtC7bDESSkSI4Gn0NXxYOdpTorDGfx7gM+63/kZUFX7Ix4ZYkmt8t6kGKgLHvrxee
/PJQPoNaJ55jtv/OC4vnU/9roa6AVhAmsJ+l1aRbEfY8o75ZpZOWAMMlhJ9Ka5kQ4so+ZFYSZLOn
73eG3fmtFTfj/yJs7Yfpc08tK35emuSuXCE6DvqW9MGodgexVnr3gXG5J6OlOc1M/y2JslMnCt3s
2EiW74wGY5Bj2MxLkM8iO/lywpRtZnrRcKG6F4Lgzvy8ZMa0ea67DMTQ7qxrWudcCJfN2mTl7K21
GywBQ1Hp5qqL9Nuhlr2wD2Dymb2F2K9rKKwXArpwnCT0ODGnM8HqB2q3Efx+PC4T2vBIc4dXfO4C
sAX2ys/fGYoJ++FhxOh8tZGp/vlpoqwBayo6pUsQFjduCDe+BPpz48kmyEz9SvvE4L7Buh7Mmj+d
LWUsmHdWD3trjHo70WngwRZUtS+aRLznwwg7BeucnTX8wVo5jRW3/vgtVU81al0poz2IoM1xA10I
Nvmg+g4c2ou2BPHBM4vokIYPrC2QU1Z80lvNtQ5wXW30/jECLRanzuRrarCtyov+Rft61/vqNDN8
2OVlxwDsUCubQuvnxLVKxVcoUGyEScsMNtnZDj1YLZQav/8/k46KV6fmRRBW9c+r5sDhWvZyxXtO
G2TjW/ulXgI7Ft91F/2SeBBONCvSCbwQ9EHDSjedrgP5d3u+AOvrO+JcBOTkuWbXLvP0VlA8G4UQ
t4Jyb5ar21rE876/b4ZeCMQiMc7X+hs8et5OCClOeWUbemOurM1jvmTY2E9zOKA8u/R9FAWXRHlr
gMZpN27v3sByWCJIQoKOCoLbPKPW2RnYNSROiP/KFih723clzuoNPhBA20Vn9uJ0HL6W4nZaZHZs
dg/GvN6GGfeES7OGDKGTBbxtij1NGrzuov/nWqPnblH2QcqkSaQZSwAb5Q6LQklg83AEa9oeY+6m
UrD2SYmXs9V0M7OUKsdKgvSo92CyIOyyDfjPVCXfg5T2rtpF0TVwnmJi+khiH87MbVQAmGb2Ymzi
qzD1lyNOmch9t+r6M0Qr0G7NPDWt8sdscsI7ym0lG0N7N3E6Swo0y/CRQVV7UlBX9/dZiMwzrxVy
JpuTot3eQzWMHxHyg/MtWMq/IODd9KGdjTfKfRAgdi+Om9qXi/aeJyYB8xfPxqmvXbzDRrFiZnJT
TQrnSK07tvn7sU4yfd3Fe7fCCgxsnHAdKZMcy0Pkrfx2SCJy7rHBhthn7xYHcLJ5mroBQlyLgb1R
3l0qA13VSyio3JfER7FTvyVF8nAqudv+bGHIOpawCnOLwsE/luwvzEXFK9L664zks+zwmBxys31W
f6GhkoKxwebcqaRz2hh3IKnKDZPN/TiJCxuyJmEJYux9n3gNUtDjOB0YC3ZxaiR/0Kb+O5kTGv+s
oASBFQ4DG35+y/jtivJz3c79MUyj6KlneUpI/EvjzCqoj0xrJWD/40uaH2r0FzL13oOSK5O3KDSN
8rmyaGB/MImB2HpxTiXz0d4qfzEdh8n6Pp1u09xlsqNGGTcf4Y0hUpMCqB1aUkGJDWQc1yJ+iMdl
8sHuFUAJY/cM/qAJFyAa5W2RfuD0Mt2NXShmnbYovODSsgTZpY1Q3KRkBjSSHiaqVxZJYtiKoses
O4Ek3Hn76o29LB79HLJp2xgueGc/bbOzpMwxKJ3+xG/pyRz956BhQRxHH3LGi/6z3LhnUGhLBTmn
Xt5Tao78y3sPqZN5RhAqFBwguLATE6S5qNQSbsp272RgBIhormvC9rQMtSd18+ZjZa/i8RG6ORDW
K+nbaUAAjpjgo2xg6pXJzVK4pkZO5uR7V9OUqNqe2dBNkbKNVNjwk57m//zwNoOffobtEALvsCaq
JADxvLJmSO5kVUhs/9jGqbwd8Yme/1AStNOlBeGEU3vkTu0kvMBACYYjZ3agcje53hpSXfJwjoAN
V/FMYpKV/lcr3h6DW4PP3XD2PWklnxZ+HrEty5R/8uGuOu5f7mSlG/PPtRFcwTjoeYfd5CgMOd7m
cuqhqXVI18O6PK3a4aM1lavzrYvn6f+Cx346HCKjvq2q/peCBh66YPQ5z2Ukh+jOg/iLlOVWILN2
CDJN6aaHbfSCd7l9PHfHirdZGk5LpK+/bRalSbLA6fp1AjZg3blffWmGsVLtjyiRkiFo7beztb9p
nj1lUZQ1aEh7xCYV8sSpnoJg6OzK8CBlo6OID3RFio/v+GkKrKGuGIkhMM8CtI6sLgXhbPaoFdYJ
NJD7PCZ4Q3KcqtQkG0G1OVMRSFrNBAPEjwYZ4aPWTNvKf7sONYS1VmAa7BmvZEBw/w374j3gCEQ5
9hqGd7U28rnQWJwgNCiTFO7Lxncoq5hi1w4E7dOj0w/kjjbg6Ey7CL1iygd6ubqfE4bHAdtrTP+6
XxYM2akLOJWrB7JPYSl3AhjAdA3/XF9TP6KYz+nu7cTfDqOb4bpCm3x6ycompmbpZ4m87pmM0i1V
pi06teCN3lu+VSX9fSmZgYlflXKy7oDtgZAcHSVvWRRrynDaTLquR9FBSoHCwjV++GKTkDq5GNcS
USmGCBQ2fzQhjkCqTTj5Cz+MNhclWr7i8g1sgKWL1+Q0gF+51axUJGSBzwP6fHnFIKbL1BUvHymh
l4e466O/0i7MiEnpYWCKac1dcogGoOfbTK1qPf1fWgqvaiQagzYro/MVYQ8daV2VOQUutnwkJ49Y
R2ccdCVlWMp1T67amfi8e3IO99zuPakucPj80tfxZH7b54Imxi2TkMD0ZGBvyLV8We5LWvbwOr3r
cfgPo/KrghjCz9iEBBqianLkkQvtruwiENlP8ZJ2MSQtTrEEpE6HGfAi2wqu7JnpoZjekdqHdYHL
QBD8lPp8zK6iytv/evHKslIVGb6vSHgA53OA0T+KaEc7JIMxyu/YLBZehGWy23ZivDoUA5Gh460g
IuFP0lFsP+FXpFecBgArZhQ1aG/0n9+klqoW8jyMCHCjNuu/blQqibTMGEQtDIkUfLd2pn/0cxDw
4+t2/zsMJwYlPw0aPc/HbCNed4EtYkeAXPZBUcO3BUOn+SmFCl4cPwq+ppPcNeohinJBcIBeCKFH
2mmHsRUEW+70iG1Bgq+R4yqXv8qXC0asrkTW0gmv4LxDEkW/DpUJxIyHWJ3asE/pb1iuVLy4hFSN
W0qFkJz80MrO6/R8ERC7FPLms7gfiFRMaWODQjR2EqG0/LcRzXm+O38CTMCFIpmRjaMf08bzXfeF
ld2HR0zjOClPMbpMBsN9d+9EcZKvo8hpCZZ4Iiilk2ItnrhuHQ3rXg4rvb7vw9EjZBm/NlKIOXrp
Y3viAMW6w5qUh78bqW2j5Y01erUrG88xXMW8YuBFgcUAVQZ1JqtPaaxYW0Vit1jj2TnBUQX/ugCC
NRTLbSUNSe/YYBlJkDee4QLmqS9ETQCikwWyTtjr3tYI1hU68h77dHsEqYQb7RbHKlVhKvnv/FOa
sYiK92AUagLAC59ePDi0N0zrMP9B922MGxeKSHT19v2XEwRhl/2j+MWQzLyHfDac0RhGIRscsejf
7Ldv6wY9owT/0mfh027D4YWbUmy3ykfWOCsy15AGBTuwGYPyuvi+KVyHuK6qa7rhopbTLQ8+1EbW
mIBWpGfRwGEy0Tvs7ngkQnhH4Aca+gJSK3DyBfJkI1mIAyZuPuJHfJqU8TGkv9ra5NfYG0As0YGo
KznfVcGGVNSkkgUt8e192qWIEh18NKFcegevasiEqlO0wbDuDd4yf4Fwj6aPeU0DdpIKVllzU/ZE
VjiOSp+EyM4bw0laXJXKpcPfqQsOwvmyyDjsZAPO7l7EwO0xH+GRV1D6e9p22U09lQP35kr7zaE/
XhZJtZMmETsy61kwm6woLZtBFxtMKA23Ofs9xjCIxkTgCJxiVqmdgia641JIA/RS0TTvza1ZEZI9
QXypEqjWgQayU301ZuOu3ClIOchpoS0D/zrPH8WeprkhzsSOWS/j2dKTnUHOceTxCwOfu3GgQjv+
ANFQFUU/R0WAvW3Qiu7HpzHUpQLmkDBS3XuCVXvlAxYjvPBCaNRGopRH5jUVFAVIBggAmne6EGpa
FI9TjgY3KJ30923K2ka3hQj7sExRrYvyzpaSo2oJAuHdwS6FmhK7wqz8Q9kLtOHugkwFLGideN+o
wS+XGw17JxmEQQfbVTzvBniWX96m7kIReZpwxk3QThYVNwVjeEOOg2eWQo6PDBWK4td1Qiq9upND
LKmG/IDZpVFkoPYkFS3xiuxVG3kEZHQ1I9URRNYcztafPVqvcSqIjGD3H6NNDPUhekwkxXwHQNnM
aDS5RGK/Ds5n62VgrcoOdsqZDzagvhQNKEf8TQzEaPavNHTVV9e6kezMr8APvgIpOGtSnqFTxGHz
dnKSLeNJUcQFU6rO2IcsC273RM00H8pzPj2RTpXCs6HURzfBl9T/lKspstGa2jsUgMshGJ9CJ5f1
XSBujwOyqjkk8l2QQfnLst7+kuHcPt82R3tDzVaMk7dWUyxUs6vIUN5NT5f97HKa9TLiYBNaFxz1
4R+aRySwYQV+EIG9rx/tdfvWUtS46x/wiqZdYyHAsLf0ifTUVjLOcEGWszNx5j7WYEG6YVak+zLA
ugTg+B8228EW2nYBiXv/ek7m2MRGXLVRuVQ7AM1IVjo3Ynk9cRbm389j7DgYvKhUQlW2IkEJ53sk
94j0A7WOvntJD1uDaHhe4qERCOuutcv0DymKXcMrP9fcQRbTRK/t0BVfpmiLteswvwEaQ7M0Bo4Y
//iN8yRMPwutKDIIEmg8UgK4rLaBP4HWZY/yoQRPFKJr6NSYlfKaX22iyrtAkFxupRXpeueDo0KV
yu51/iDakEz6YUSpUbKhUeZqyvjpSJLOWF4V6J2ZhKAOpGnKlMkC5HtT+uxjev980T3W1Cb9w3lU
rOp95kJ9i93LYPW38Me5o1zgZl+RgFAwDnGPOB5odm0BUookM9tynVVXY1cyEoZh/sJXQS4qWTl1
PvaTlTBvEjQLbyi6vN8MNtwXuzr1FUoT96zUChydpHmrlJOlJM58MWz7bBvzecFYA01NLm4uQb2o
XIlXXlzN1UY7e+oWe53AMnXAgkm22U1JVlPpOGAkBs274BLYoKufraqiv13O1ktdZUop0w8fWnV5
dkM1KQKjDfPT3RE0wtcyvSsbOF7+5dzWONpbtj93pn0D8fJujn2l91dpFRGPS9hK6TDtgJeIm1jF
zcfukcQ2e+FgLPsx4g0efVGeQzqH8UCpqPo6b4FbCFn3BslC17U4pzio0IweTXbKTdsjHnQemIYE
O60GZgfojMXthxbO8CdMI2K/mpZjATd5XC1QwV5aZnuUVvzogVCgmLH60CdgkLV6pDEBnCyLo/lb
l7gtXikIqufL93aLEjdJvNshFJkxa9M+729l6YuebldgwRM11pb5eobhXRUet6TXyPovIlh7eQPj
1eCZM6ARGM0IZsBE9AJkzDntwEYtZwPOlnF5HmxA8TL34vwF73hq0yqCrDAEg953JPJ4M6ntro71
yoHYbW0dELH/MyPzqMOo1vDrqo2zUp3otbIEEE4wZIPWxrZClkPnBvTPoHrcs15jLl+Bydut9oZy
hNl21lJcID3UqHJ+WWrWPPLEflJDS6CoTNVjSkcMf1IEj45axo++u+rWBGhHBmwl1KoUDdU0srR0
7VNZW/YcCqfgDB1dC50LPedoSkebHHxdx8Fcveg5ZVuvlCqJRQJ03cBtwAQDzn3ZCIhrCyYCIc0m
un/JR4ji3mXf/BNieLx07zvj/YTw4fdl4vSpCtn1jU1WXWh+G1JjtUfDc1pmHzRTEOFUO6kwvEQh
dVVAT+mDSusfvX3aVF+a1r2H5B5+UNqIiY9/GZxbTiwLQMoMZuQOdvzZrh2qoTl1vpBlq0Kj0a1E
Psh1XvpubFdGzCA+j/Dek1qNjF2kpe/KYxZ4NAvDmbqgYm4KmicqHv9XhChwQEVrxeIHaKwGJyIC
SVP1B/OHXyyxA2Rny60i/uXxI5n7MALUvgPrlGBHcuVWE1xzTVTKi1Ajk2jL0GPSjxF2vteWcd4G
rua3vTFtRvJgo97APVpt/Id3cmOGZyLx9BEucmkZz8PO0z6WCrjo/SD4ULUWfb0KZnCTBSOMwwuV
IH04h+08FnKbtSSu57CW8MLekOOA+nPsN/rXQ7QGY5arymgbOx/M/jd4cLB7SUMWoTRA3FJrvqzp
pj2obDEzfZ/eDhTPKkSLXOWvRO2LcKMmGpMSURBqAPBtKNFu/2WW4k8DOxxUfbyFQY9ADbsvh56L
0RuaOGcnR7ybF7iM7FEA7CFo5pzfHDrRHP7RRujDzIsiMpygTTj3C4mfGkTuJjMhkBo2j+AeKjA9
k2jkrg/Tw+pOQEKiOyeN4EjttbqZwaYUFd3zyErxRCsCTK+dnm1Him3f0MkfnrxKAON6VV8OwQ7w
eMANLbLCxzcizQuqejTc03fEcILuJhRx09q1XgsE0RU1ggEtnaOpiPYJ0k4GvBzoirTdH+674vDl
eAauSeeNge1eIHbIW6GAu5F/PU/tWsMbpcQFmaespveZCV1NfuZ9o5ihDP677QxxSYIdWA+wBWFU
z/iN4AAMG30iSZrJ8S9i6qd9HN8W6hU76NIPA5n/9kcQSKv3yN8Xltd2USEyY/YsLTpSatd2hB8Y
PXVgasOmWQLEEZ5X4eTKeIOVWhbd+z6Fjc+T4RJDZAASw0ZK8kSz8zdXEGmRLBjl1YSGiZcjaEU0
NWf67gBW588GzcHfgEMBd/UACJ9pf23hVznTwEZdICGV+FCjkVLYp1lYva3y8snnIhNKPLg/yAV8
7y9Pq9AQfeDOjxU6c+jni/gaZEdunq7m8lHelUf8hjfVUdBFoqqZUe7hzdb/4MTN4zYEHeLmtr4t
ndWv+saR7wy3JKJKoMm/UrdcviV/fnSL7t+Zk1A9LicGbZdPInec/ef9qKdTwbM9Bc/ruiNt5nyy
kmlOzwQzhkqaB1ULi0eIP5NTmW1Y9gsVOROw8R62a2bxZouJGwtpUkk+7NofmVd0v+s706mWYKw0
yTNJsKpDrhl//So79fh10NMCe2k9QtBCT5QGBjd37y+0zH3aJsgaxerRCuRRHZPvrsyywtbzb6QA
By35LtuxptSKlzdX3ufh58CY5BHc8hZEFI8RDlAIo/Kmh3LZdWUcTx6Z8xXll+V6cRpNAiBStq/I
cD45VSw5H0njc+1tiB/Wj2KNCDDIM3CGlMYehm7m62pXm5UCbMjruhgW7aHBs6nOYesrbS3wfJ1b
GDrurwgZ7m+gkBEcs++dHudRLYw6a158o55w4g5W5B+F+RLpNvmvq1i9gecj24CIdnHkOJh3vvei
8SYn9ziHlnPKTcl1TPz2wb45lzWkOxKqo38l1FPby39e1BQWwjouBoYtPNW7dSr3K+w8FK74FG5d
CkZnW7jbnbkTQ4/KRz8emFgO45hgJcaZp/ChY2D7mZrygN6o654vdcZuPh6RcRpz/e/9qw5IoDvv
F4fKH8BvOvTybukr25I9VcJolP8P7EZQ+0nmW1Goz2GC3ww4Pr44GFpaEuVn5BovrnAzcgvME1td
MWF6hm4+Qi3XmCBoWVeD/PW5x7o7gEXC/vVqYACwy6hI+ipcHsEvrHtU+QM9geduJx/46Va+f1fi
/8ZK6PYWD5ndfRMQzpTRnJvpe+BT+Yn8T1V1qCoSJbk+62lcM1yMt8x5TZye6SKoHKJaGHvyhkWs
s61tWEQenOxSQZiemoRLAdGn7+aR2cINcUSh0z4qClgaJop9PDSKGmeyZI42xMhHBkWyAzwiMWqY
E1Xb79QVGKYhUcRTfG/eiGIINiqn+nbMhAknmnE8Za2fe26VEaV0UsLLou1bUppnP8kiEHS5EED3
oaf/JfgM3cKLgtRuPJnWVENYj1mlMy1aIoe98+P210l+/6cHPO8y0/T589P2jbR0BmJTenEFjCpS
OOKH9H3CvQ9prpwoEmJfpTF44oZEtG/mVpR6pRiK4VQgQpd+iMNfMYdYQpkgTSPSaPvnzxMuZakm
c8Qdv4CfzvdZqD/BzRNQ3IsSilHDisi9vxalVrU09n7ZJdyCHAirrMeMNb2JD9GpYG5WnLIGU0VR
/V6HP4hZDnEx/88JulMy80fvtUEV4db8dcoJqf5r1e3os/9+SIW/OKTsOB45XPptGHftFZ64UDbB
XKCxj3K2vfuLyho50ucDhbA0RGdzk7mbR/OQbuRs4h0gK6WIBq2akqnBBngipX7hH9ZShkfpLnpN
YyxZrF+bJlRvWni+ujSwYbv5OSO59aPyVLvWStS1U91WSIUt/YLDxT4q+gfECawN/+OjByYFU+W2
4AQZyp2baSDCq2fj77UUlhKwgl5c04PzY6b04SHUG5R0ww9F0MtV9fd4VP5SUmrylD3kYgkwdzch
9MSYDpjW8+jaRzZhT7BHzlJP+kH9xq9Fg2psWRt7Ufz1GEUo/stYgFUKafD3slBvEPhwgXeDMC4L
eUNqWvJVWXv0TikOj8bV3U8EKIRrBAI3tbq513lZ2XqFci+CXoIj729GKURCR6v2rGTVw54Cz2J1
AaVI2q5q4Q7IdtNAezK8GcbQTOUPElfbpnZvi708pb8Lsgm0Bls12kVjsWSOJKpUdpvFuZYy5hli
gctpFjZ9gImL7hJo3fGdVjfMRlVnamVlMZhe6a8+kE6fleQJu0274ANfHjILWzwnqlwmyjgRJhaX
sHsfIn/DNan9waF5+DD6H5jffJcI/PW4NC4g9ZK5D1zjeFeLaw/tzrQu5cvy6HkgAzG/GaUrvHRX
GwMjHqxVc794hQF05T0hncufhkyP+F7HVQTYqyvmVqWYsgJtyVt1FYkE5wNhE/E9zrPhrwQkHpqC
AWW6ojX3FUls00jJy3vSV5iGtgIf0xGWtcEpAbl1qp4oJE7FvXTotCaTYpjHQfK/lAdw/no7y+WU
1NxsOFGBN2hVdZc93KtQYUsATG77S9hHy35xlJ27m1q98cjN7m9b003PNbGNW3GDywn3dxr9PTsA
ZBAMiqDWhunUdjopnGr4I19nV+iMTnTRSJOZg6nrOAsjSU63eRnvjgKX8kM4rI0qkigHv7fVzQU0
dIYCm7ISsXstQLSuNp9Zq/a7EM5QXCU2TIuBRWKZmcSwwszsYabfhw8bw+TuDIwTsCXkXTX0WuLe
2PCi5CvUMWem3/nxz5ObG76guunZY8qKCYqsrM/nB0tzhxtuQJn+S50ObjIyuSjCxWgS/lIMlhaZ
QXFcM679geTuHDgf1ku1plnhu7wuhV5mKSbksSQLyu1sI8FANOOSUMKNbLQNeZNRs3TM0BMdVvFu
pmSLe0XyTzaw0tjuNOC8jyv+H8EBN0XoML7jRXvmPXL3ypp2sS0dqIaBVBdlVIhldpk5M4zr0GKf
sJEFDUegGeInbIbkwVg1xSW6GLbvCL0EsZWKcj0pDQihVxWCBI0+/v85NPf06WjD3I6Cs7mNczfH
gNil/V5so67EbRMxWXNDtk0si/ma8K1Ny7pnV5Cb4hZPYyfxVu/LHdOTxBwa6kDJjYCh82T0Z3VG
ZQXS/QKNWrrSXibXLkh0cu5eHbewWaGNOF/k4g3Sexwa1u26sZf5ps/vnrtD07CIIsQXyIkAYSYa
rGFpv6MIqEPoL9t+SbvVbmvUNrGLihbsRRsfU4OzbsbXFJbslyxAeCtYqJBU+7bPi2FhW5FWPLj7
CX6GvMmEvHW8W057vvg7jLt+UGYfp5eHxmV9xL1czcuuQloNALcv8MylP4//Q8lQI7XdPGn8sy3/
MMPw1UZqd/0ZTPcWuKxKcHekzCzFhAhBbtJNncFIrwzBrNDBT7FPrLOjnnv/eECTe0jAs87xap52
wHzOHtCnhKhmI0uA/TifpfnfIX9Z6N4lNqkV4/K0GNuSEjpOLhy4/yJgzxJF67u/sDAHQzSnweYr
9NyVVQ+tHtxmQaZy1mXPZuHUKNFzqDyUA6oI1YHFD0sj1xH8V2P9KKy+xNW/DIpYy+3PRNd5q+vW
N50YyDeNkTSD6P5AOY1A/uRK/ResTXrmdgjyhkHfbPQqL1dmvT4I1z8TTiAOBQKpy31gG0P0955J
JdjDKL02SIUemMvT9kp5HUaIuG0IdxDSJkycTKO+mJoG3If/GiRv56xEsg+JXsAnfbHFExUzYm8i
X/k8jr2zYpzTZeDcN/kWS9w6TUwodDKacUfR3I7XA/Aw6WbbED9aANLdkRxU3RuSAa+VKN7+3RrP
FEqMVDNQI1Xuu/XzCLL7bNQ8HqUbvK4AdMFmVXVTdUAhcUw6V40XN4heEh0v7r0jnuJ8vkbczVBF
pdMASPM9aff4g4NoOhQwC73vQ6MAoh2MEZ0wEvpX0mXAdWZtZImAVzFrvS0NMqx/A/wv0rTS4EX7
I5dVc1YuGiqtWHjjeESQ5VOKgarRVPFZ3jShT3Jpsu31SrPTpLsVTEEMKaQR5EhlD1/i0AkhbjDM
KJooIzEyCPamAVRhNQU2ZEjioWJfWMgBdXdZkN4Njq2sJ8oCBU5XCKbl9c3XnE9ltsPbJoXSQnLT
v/5dsQVIbJNP4nyk3jCPq6jTr1TRMQQRX/sVTrGPMR0Dh0upT3CyrKKj9hL9RfLVqca4PT8pAAP0
YMBzaDNfuQzVcA2mGLatBuGWNlG3ZjxT0jm/crvn34yvVPs+b+XZhomwOXw84Mq5ZVZvyGRJT+Nx
QpwvtREMgd6D/+b1qbmUoAtd43wFtc8zRtFwA48hx9KCbB4YCPBDOwzJuh16Y2qJn9Tkc5vpnrbw
mt9A09rrxtUJVbv7I3pJba+ME73b5GogfrLiLxAaYLaYk6U9w7MfF0xpQd9Rfb9mnpRWeo57BX5s
T/ajdtf7rvzya19pXA7ABAMGw2B7pZh055wq8Z6jZP1x6uQu7w+KoTwE/KgAVbIRb3DdkkCfbXs+
zAORNh0r1GH/ZLeoyv1gzQdy8i0Secnwp7nB8MXR3YtAD4Eri3ZkzAs8COqhnr8WsHbmvjCu7FoU
S236HqmmFTmuDTA/Sk+RKOys70F1PyxpnVz/KBtjN3QxyD9pWii95LPfLMjVY5KuEkoD3HdL4ZZC
p4jZOBR9Q/fn7u8tWHH5ILsrbu4U6lDzJnnW4cQayygFCRD1jJXrQzaTndUghVxnb3qK4KDjMvgH
fUV2BZnQQc8OoQoeG3r/em1vZP0fjcVGSQTBSVZr5nkvf3BPLFo6mHhr2xWnyIM0ro3UOL0IvSne
fG8cwbuz2GUrPdA/nv4J6zt7fIvl7WfT18LnSMbG+zTH1dqZ4GsNo0dQfa7E6vlEXDQLI+rDoJY6
Bnaryj03txhMWnPfyBPejlvY0kgUXr9dGvok+Z7C7TYzwcDgFaF4SvK94lUnnGu62o1Sp+SUIDmk
/zGw+4IJigVhxhDy8MZofbPY/nf8OagLS5cpdkzbjuBkAt6VnHLcYgih3KKdNjf/K56n28TfjOgp
1DldvsHEzNflfBSEzOQhJYn6y7AybNRDtcAAd62EPJ3wDfAWKQW5FELFpO9shrVLMoaziYNHTXzX
1E7USCMbu/n1fmR/rkOhSY4yBAhKyfjqyoZkobpK2i+Xa/5PkwkM6IElRUmqYsKdmN5390n1cc1R
Ed+JlQDcKgwlg42EA/ulqA3z94U4RxkjXgfOzUXYf9d+XmS4Amij5SUtnKCw124XqGqKhkkB2Rbe
mZ/xPfFLH9dyxAy+oIgdZt/ouBihnRaKvl/zU8k/erZdgIPnN3vhQSPGl5qb9KJeyB9I51mf+OeW
L6Hri9WrKmIVF2rQ0WGJG3xbeCFVsjsdW6qGlLE3AmjUCYVD0FjSfQVDrPficveVGkX5f+1uESn8
LLczEV0V7vPXZKxMv+F01/FFVPvDQJA1RBZwDNDSOGaUv0rMG/hU2s9z/1bEEDd3nf2Z5DEeOe7/
1P9cT7bh8HxcHq8WVJ+gKICKvIpNBhjOYd9Ebg9i8TZf9AtNtFUVEjyu8YXbLJi4FgpaCHmLkWWI
GP8kRxreArWu2TvF5JOWIfXyWDmYT3DFOqdilaLJF+pfRCkHnBWa7kydbdGLzc3oyE/A5Bp4FHgi
U4McWH4xW+yjy+4Zd+zPKsNxO43Rom31spC3Q/va87PSwobaKH5HX0kWC6zB+oT3rZD4eYnLYhAy
5J1wEvP0y1Cszyo9eC40Wy5ybxVTTjxiPDyNaNc08Yb052bWJGkMCAtNdfQI3Zc+4bGBdwDMp8u0
OiVnR3AiQAIbthapwEoZ+pVI+5EqS1tuhOM4z7TfjpFisrQMbngYyVnavtYq7snw8WBwfNOO+eLo
UUTPOB9mq9T1dBe6qI5GkiJ688L+tzlLQnpcLiPvaCjTdkicecMzkaML+HzN+e3XmP7EcsTBwksJ
FZUbYJBnjbQjG0rvGTMczvCeYYN+AYlctl8Qy0fEaP6JV4IUSJGtYLdM2wZx04ciIW5k1Z6rX3vm
vXmM3yGjbarVWJ8Se+sSRccQpsX4CF+9hev2nNZ5kOiJLLyX3ubfzDbaAX0MbxZKYdG3jlul6EiN
55854BqwqFQ5PdOnW+XJ0pl4nVpWEu88AbkljlSiKqgG1ojsSw8hfytWD2KUpExmUQzYBN62KROk
mX7bGrh7z2Kk6Ozc7mfrAi7I2VtBVBJlAeDSYRs0xhNhZNdvqzw+L9SWl/oZu3OpC4etHHkOzryq
G0pPRt4YbqPf62/XZpGJBuPbtduYjHQR6cPTOIUrvFOlRhlQlE9ywU3qtOEmItHjn/gU9OUKuSEQ
dw/f8JLqZrzYK1+Jd07Uza6O8P8xNOSOAUUvqx/0WE85jiOEg3HY3tElewjaD/FQxVVFDDwnGdlR
eLGeZywifyU91HSAArhUpO1z4Sovs+wwHkJ6iBYeoL3JGA3tsxE/CgPMCeahlmInnYBjzZkSFNhn
Lv6yrY3fn16lnGNlkHTDN0G13HWe6yrkOwJzdMtw4aekozYuAAdVIz1tf4IObIJZKptUnZg2oOZc
r5jOgD0aG9GQCpAPjAh//zRQ+PGOxksqkGqtS14R7HLF5PaGaQYqxB0mgtiEd/TVQ34SnsSJ25ML
vDO/TyYkE4TzXhxnUTzB1CyQAa0UBLxHv5vwBJQUX2OMo1VFoWm+Nx6H8rh6h+AG7K1rt106LpDD
e14uBB/RCn9c3gG+/DmTWH5uTv7rzgLz0m4GH+0MZAeaRTTevb7ys3fqWlBUfFFijAG9EfQ1yEtN
RNNvAQcHWBMyQW+lDg1Sl5aPZzhVm2H58QutgZBa0HZdU8B2DQ1tqsfAVT4tKwpdzFBRshdtSSQl
Rf66KErbi1+SnGLF90e0wqXFiZ5jcikl2gJ83Gb6WDe3HJzwYBOi6oKPDQtl20b28jbq6t/bCFc0
yL2EDJwEcNcdg2RbvTeMdOv+FidfGHvihyYuby1o9RgKynDg6/BIHlSvBHIsAlgLe/K2QryugDZd
LDNzYSxY6W5j4GA+5+xHQJhsh/3OSW9fmjoiNZJ6NikyB3gGBP0nTR74hlLQD4+J0IUH1Sjr2RYK
y35C98u+94Bi5L6ctMhf8jvWGI249ulaJQ4JmMeCTtV33AxoYg90fBTXxfjy2lAUdEoqLSFTUK+e
HcsGGlhMR8j84kZ4zkFawCs2/PVFPNTYo+Q8mSonzaWBTBf7tj9J+YMmFl0tgIJfatJTZfYT9meZ
eLpyqfiwNEMPmgDt9pFODMb9ZEmOXgbLkm0q3cCl4UZHf8Qlckb9BRO5RrUlqzVh9xHwpfEJU7Cs
aHwOUEOqWYLV/zUeCg/Wdw0SBlUBKYhjRIiCoSnd4Z2OY5iGgKmECHEoAR0fDyyXocN0oX3QbMRf
yW+TIy94fuEHzEDUyaZkafy8kOlG2vkea2fzfBJ2UFPyTbM3PwqtHrfzONvEQP6qZVDMRbPczW/Q
nT7q0pRzKUKSlMRvKqTxJxmv+74/hZ9n1LW1cP2PwjEpxYWhBwDbpKPjG3pdQtUYai7vAnIOjKMH
pPNBIVrh7b+7+JeNCfgzmfmgXmu4F/IlCX06oGRvA5s373SH7Yj4XxWmzWTCZeKuLmIVohcIlhcX
ALaywAEEpuzyUau5YmRWSRJcpiVXRTNAcoFaOikwx+zTcTdt4+vrCyaYT/IeRV/ENjzVkI1h6r6h
F78dl4xFCf1VC4hU64MkpNqWPRexQH9gaJRLve5UDee8C2SBK+6YODxI4FehfxyImTJg/fW9oVXo
vyXpFxxMGIjlafjHh/bge6PkTuuFkZ7XwdiJLl/A0/EbQgxBxrr6PtES+8VMDhQFtA56vend6nJZ
gJ4C8SQ0SINICO6FaQDya+Zzez1d8dECpe6+HIucgWBXP8f+mFP+/wfzzqgkM+pRRsk0nAkTtPnq
fjJYsKe2COlImZdu4SbNgLpnUf3LAgEXh5zO2z7k7E5iduF0AJjCvgbTXosvZTqBxnM+qswHJIfS
bIlXkPTCaGZX8R33/m0/8HzUTSibzT8joqdAcSEMwgxTWzKBA5L6BzEwXCqolfaIhMIZYaHLXio6
V7cMnzt/YmPVaIUFt47EoD3zFPUJQZsiVwOTjFMe4XQxlzQWd0aUQRiyAK/J71tedCY/cvKOSlC+
tcXgh4gILzbjf03tEUT6N0a5dLFfEyO7fgyRGF5i0Dr7cTGJWKugsz1Wo5kTyYsr1jKfKrmWD5Uw
ABZUuKxFv4FW5QiJ35/ksNPXq1TyU9wxl+/Z8wD5woDO3SHRuYpCq4RV2Pn01eGQHuzvwpbWi1qH
KvoFz6qjCFZ08GEzTm+V3ExWdXq1tCfjoTY9sHdmRyRzwgIrYYG3CNSf/SgkY4YOiWNjIqif3eXc
Tz68paxFMTEcCnjWOseE87d5EYYggz75tC+vxe3FCo6+OnN7Eu/82XPJrO7UJC0mczO05AbvareA
rjG1sy0r8a8jqURor0WwgOzff5huzaX9FZHCyodIpWa/+OHBQbaEpB1YnAIo1bQt5tuG/IK3OYmk
ceN6X3z0LcNIw2OwBDGWHcra2oWQ6JWoaNa3zJ0ZwcJmYFQjhomv5p3Ds5RTrNtIc+p2Z9sPhd2j
Ce1k9MQTZrPQT5wfOI5nUvCEvEq2wadTsoER5Z50HkOniq1A2mlETL+k9tsQkvrcdqWVxVOJTX5j
K7iuVTW1btFZl3AFUxEdj9vSfLLgRsmLCHzCg4Uo65/DusQAJCthhTyxedDDeQ9MLkNU/LBSpjHl
PHaj2Ji/7mF9RJezPsCX12ykL26XrvtHWas6URIFy+Jjgqn3Q0Ud2p0YBBnlQ8LO5vgA1uZ1Wc3k
9jP2Pa2ZK7wffzoFBIZOFsJX2KJ9pX8bNxu0HrDLlw3nFkNgEVFcFyFQV/whN8NIo0SRJT9t4Ity
O2nQACwZXzqTSTZWPc3JjinniqlxxZ6kI2UWo+SZ69Fjff57gbId8htEeNqRTGy4Icl32+U6Tw8X
gAm6vWZKuU8Q1AwXCVUaflmQGPMtBjoo9r318cqXyJalYJJ0M030cqas+38RWHe5wQiXJq4VXXdb
yhcMGpXZk6KaYWcAMgH0ZOoV2HOoT07YcgPTQHQWBcybL+ukKUARn4WMROtofTNBSDuNR1RPah/8
cql5FYtOlTYVRDEXLXu5S2zq/FR8DnQpJ2zHAidjupEiTXAW3m8KcrKQsd9OnVLLKGYLhAlqd+WF
GFS6SNuAmimFxTLqHLnEzbd78m2FMaOQbuWBgorImx+bl/IEtgEiZ+k8QSJ/DdCRjCbbXJDAX0He
4QXhUDICqmrjywyfOljMlOiPll8kJeO8KSUNizJFd917ICFe2qNIMOds2GwX1HDk3UDAfXTfrrCo
zrdLuCNZbtnAAsSd8tvSpz5LYL6WN/HZ6Qyt4qQbwV6ZkVlO6SqJM32+pght7x2xfq56sUE8snb2
QooP0cR55KkwWsNXLg7TjXxDj+UganVUCAgNEXUhmeMIyBamSuhu9xrKodiQbxapYDh5PDuNgd4i
5cDemRQ+NtnOKXGvfE6HoNOzvc0FeYOOo1EXc2P5Q4QNsQTCW2qY7Mn58sUS8FoDCy9u/Ruwo7RJ
p1sCzn2wA1t49WZD5GeaCb3PWTFuniuiJgKKXci/k5WE7KkdqEuq5iE+skvDcWCbylTJB3BY2kJP
T97NacoUiO4Zhl6g6B9zxgirN6agudku620Wrv1mgl6mT8c/qh2Veuwlsc84uUJf+KnvGEI6B2d2
7Grm1ZDfpNFe/O+7hTS91bfDpC8F0+jA1gReN+h2hmiQ6f1IjTkuw+Gy/G7RvqHp+UXLzcyS98Zy
cDQx1o+qld68sj+V8X69sfw1YCqqFVwT4W9uPm256qmak+c5qDlQXK+JKkxAuun4Bke4Cyelrh7u
GCI98xboRyWMd7Ld7Xg2AimDlu7OgVEWQnXGSmpvgBc3bXAOy+7jn4EuWJ8gG5L0FnqX7vvlYP6s
VDR+07jNP8o0i2oLQ0A5yxtTK5Aa4oYC8xZOhrEaGSMtUknrjZwjKkqp6RQJ6i8j16c9jISdjv+B
Gjg/FuxGGmYsYazdBVhfTVm47OagV2ccJfmHqa9uQaOedhn8v3yAGQDAzUnPWMA+MUuPnBnY2XAg
X9S1gyxZW3Jl4hYYN3TuPSNkAqT4OE+c/bqMVtYEgsHIs5VRuYx4a8VB51rvy24e6+FRoM2Ks0fG
8lCzalUyDVsgHDTPvUlu5P//2kmMVIoshsoNy/gV3s+aSJFN/AxLNgAx2dIp81ovSSmPAuudceBx
Gm3kB1EH4fVv87fRGQLmVAzoUFUEqSQNxWOLAgFHdDu/ZyzK30q0a/rThQR8THn/0nHwoyRq7OJz
JX2CQ5ivZdAFh0mHHAGVV1JvzBcxvwLJssgELNH3x3zWmCl3CIjY3o3BbluWSS906gfiF4ez0C1C
wPPy9UihCnCtrKD0z4Ov6y4gJnlatrDdBdwIYXE14a2xPuCom5o3Z4BPlhfEweFlMFzrWgan3xZt
E3DVVDrZUzYXXbrANnF9deTi6WS13roWUfkeU3WVkgLt4+pqINvDMbO4uPqKvxZOfQC5POcZRRt0
H18EAxcjwqpHFJ681YeD02fztMAFLkdTJWVJRiew8K/12MXTwFWypBA4I7WnhDoMdiXRuXgOM89O
1Fj1ueIZQi6Weg1JrECvlIxz4cs1QpecP3dw4mjQSzcm+z3l0rxbZy0VDqF8fvbUruDFsqkmRKsS
PGUNLHU+b9wTqvN0hMYWRiamMS2DIA0B5BAlYEMa1cnbd1tVhN3uulx6mvEvfWtWwFxa0yWhii39
6dhi515KzW6BqEtnRnun/Us9uQroxJ4CzgkhzAAVNWYcKcJBtb2LbTaZeL+Hy2xHSIz1MBdZhdsv
UhD3ETFRz0M/aKnn7TJb361LFIs18MOd76KuU7/6KRg0+aJmF8P4wt7L5CEvCoCnRN+ggzLDRKpz
ge98Io653SVDnHmXPrU+eXVwKcioK/dEv6OjxHd8EEzRRq37JJ1fUhZ8JH8bCqxjtXzB72NI30jV
2j280gNbvzWUZe85GXuIBKXr6zO7G0f85Buij9EFn9rD0A8ma7Chd6LIph31LqnIpXqWbYXPIsVg
j9Ag+PtbtJ4e3vwOefAKLXpoxPujmYxjroyw6QOh8P2n9PddEOOnpaYuxGSGKdR5P/PHi5o9Eg3Q
JpFPVZUbeSVHOKWGinTfPNcCB3RTwolW9VGsmmickVCthoh3VadNDsRcmWytrz4LfxjByP2cnmZK
t8MPWPsytAPWt4wWtQO+B93FZT7IXVxliTuOFzN90BWvg6GYYvlfj8Jhk9kTVW63GJXW0U/vTYlQ
0Mhb7DfwBwmKCfpbpOzs5IlxodNUv3bjvIcePc6XAldYR3qyGpkXM4YudnykIn5ruvRNetZKpUjx
rr3l8KYFhNNbVCcDgW8uZkpUg2eZersyE3o9kqveaeeHFU+mP7Jew37/51MfOhy4RD2B8iwOPjhH
PmBg4hgL0ek6OAtAsT6+vGqX1OBEzGJBweyvd3Rv4cy3qOKvHEmbowvV4wdqDL6SZGUZLqTrmwQS
M2/oQrAuYtKYWnp+f4LqQ0W8x7sciIVO1RMnh7WbK861B0YEIz8HkeoGyMGu91pxNMO5ip70io/E
HvLPgmBagq3ms36akBz3ilZkf4D2BTnrps9l2vUmCf9U9QWOnRpoPR/Diaq/Wk9oXUKo2UhpdunB
dhGMmztyRd/rgVmGopM/9rhrJh/yuTbHsKzA56wuVsKere4SwOkWojnYK2BHW8PtfVWx704pyaJB
Kmgp/Tj6W548U3eJMQM2EV8bOHXAj3VcJMDVCNgpGe28ZbaFqc7JXjpcx0XPYDRnLFkkV5amhd03
T9knNKM4aiRVhCqBxXTZSZxO1FRyJ9vsopSnWb1efXdOTR4ZKKo1PZv/9qOgYuV6aAPQQ5UtTgXu
bY5LMSJLDaX0nRBYXPQX2ld4QTjgLnBih7oaHdShDRqKJpLBbyaHeFW8HrD4dCteW4uGTu22VaVT
5aQdLpOhiWvmipoY9g/zAEI36dww2TqiiiWRvXuCRc4vFe28SFfDp02U5SVBTRZ0zpVAXoQFHrpf
Be8LWjOizwXXznJrUmgx+VpDSQChyV6WJbIcsPBatcRokwjIdH2dZTdIWk31GnKJb7R6O4N7hGNB
haKXF6hOU1g/Lku9WhAhauzMKCqRX87cNo7YVteh/I579dou/FGmOpmqBWFYdt4qAwNQmTIWGyOy
+5oLQgv3lRB70tdoMP3MN8/HiTfdzpSgksSaq3jkNrRb/W2B8tb1MjNrkKrvPHK/ovZ8X1pZZQfw
2Lo1ltWGxdLqAjTmP7UO6KXLVAcleGkk3HoGSf0GFa69iuHbUBgLc/1WxL+Lix6/bVh2qa4loVD/
f1GzAZlzS9r5LbBcTTbfkidM+1QsaleqjvwicTidw5O5iKxibkEB/CRXKfpjh2n8EX+ow2LumYIz
bUBXk9X1XWy4Bvp8pRUjm2LSHFANMbavhcRxQwxHAkqvp0MHB4zPZhaJ0SbbdeD5lWoPXS3vm++S
S+1hPH1A1+UquGUn81LJQ/L5DP3qqnjYNSHB/f1e30sdDzr+9FRvkog7fLbGQ/4ueFEkOD9vg8Sc
F0O6M32Q3tT0WxbMBXP/9NLiEE4TO9cPTptIgkDWNxkQoHKaXanNaZtiKPZ1fay+Hv7ufC3flcvu
UjxlANMNqYSwgDnzL10QGqibgKD57UgdgwoK0pvmYGsp2Hk8Oxie3p+G8zW3uZzCglbou8TsHtvH
kWmmyGiKCCpiMpiFZzB6neuK2PB62J+HxFc3regCj8yzHPuIo12ad/GbVfSo9Cn3iLUtN8SIW09R
6FwhfbiJ0d4LCUcPR3mfm0Ho2ZZ5cFNZfCKcntlXS7APtEWJmFmj5SgHaweRfKALcQXxnmLy7MqZ
SRp8AhCmZkU1qaVfJbw/LucoSkaqxQjn2ZjPbieuz4EEobxLSXFLNAOkSJpFhRk4vZ4XjKWkAMdl
bS/Sn6Kr4sVEfHZLwgPcg0MH4pChNY/FOVZoJfCKm7vmU2IihB18YZ5fajWOFJh2mfCg978adAbm
j1C5zqOX0gBBfNh0wUxoprv9fncDNDhqXcj6FGjbxLgnml5CxqcxTP26OudWRLalW/l3S4bVkcrv
ZBhAL5/QsmfLYTfFBvn75I4qP/5fBLkrVITZzazpSzTdbCt09s0xVEKm7xBAeWq5YIql4PtbDLO/
NoRwzOceR/hTZo57EdCV75XOC8QpVm84Nt49x3XQtN3SiIfmeTCcp9b1J9sLOTYMjI+J/Ve/G8ml
hU6O4uWi7Zgle1lNJn1Na2gXbmBim3LbFbTdKd5dPDF+aVYa1X7/FskrAGxBYJ51/nX5j7Ivi/Ho
tkv6CGfMaj9tUDknSfM5AG8Tj9J47RBFZJQ+XvPiPOsf4eQ5mOmxejkz8Cu2cH0Q8gMNAJTg6g01
nCBVs8197EGginLWpMeOCKpjCw75br9vcQMGdbEpPHfe7cfInhG3eKCPtJQNGHgfUx+jOZqmfAGm
yhK8r2wcyogAjDTRgnhIlBTo8blfEjWvVB3YUwGmmUiVt+mOex3qpn07YeNEFd/Nqvj+XFgwySCo
LYepvTjqmq08Zjv1czVuPeW4qVvy7RblruXLmmVO9AvkrunLm2WiUNCviscQ2V88WLmQ32dZIOPc
xj7Z+mOTnp+dov7y0FnCP3aYRFXcMjY0NschH+EwebqPRnjNXGUZzs1O8D8yC1bj3IBbUIdGdAMI
pI1l4usumUywnofIQJXdei+JOAwV//Nrh/bm5/l5yJIGc/URUL5qK5HV7vqhuto4ybzCzStChpGR
0CZSn0N3gd/M3X5a7ecYNfeY/o8KnvFOIVBOMHlfeeulRdTQt/z3AES7kEA7KRfmR3F+549ernWZ
QIFhh51m86o4TW1t6ovgA06pdeXLh6XSpr+Xg7lzYJ5w9y0oKN1WHtsmzA9FyloZo6vxeXpt+VLj
6xI5B7bSlZWnCyoR+aVohR7Wo1EqqyWSsq0CmUQWGdLE5yzUa/l4//6KVeF1qeVjlGgR9nzjU58O
jDDAbrzL64M6eZ1ukFnMF5IMHVIorvZurapUS8B/7hFilll5jIl+lso5cTrfXj+mDnr0LyMmtg+f
oCZGkDS6xT+0Z6/LdVoiv+IWm8XrWLQffdCJdgecYTEVibemYmy/zZ54viVt8RGbTqqDB0WLJkN5
rFq9bishx8mlbot011aGcvVUuOne/qe9CWHoM+B1WNRyjrol/r9cqLTX+Ga87NdKkX0b7CD/HUdk
+12mQv1dAvo2F/9oqDb/vmwf+yOMNHHuU48bMJxrILodOqDvcyQrQ6tqRJPHCInOkPrc/ON/+TRJ
W+9I7wI5rMZYTHy3VWAuoCDEsqQIj4ET8ea9ygFNIHynqk67EPtzWYXqtqLjDWLBa3lC+s8xiV0J
htY3tPoUmkBxY+ySfovdctImgZj7VLsDlhKIv6JNZtcDD+H8aIlMr3iSjb5VmRZHoZubGD57VEMR
qR2VHRJ7NMGsYgigQkQZyEbml7LM54CJafGiIgEjpofmzCFudpfQlopNgQDjFe3HOpH7NXgvvcJG
lgwwvBGuwhSFdR72kXdPGTLdSmQEpvDupjwevf+IXQqEn2klD/OkjWXzNLtplClAr8JF6/XlUZEO
/Eio7G8NftYL+snXAOxKr/wYXdeRd1AwIHQP92Zf2bY+fC5ig+paaUP5NhAudYgBRds0C4oSJSwR
yoNAF0n7ztUveBh30uUOUTTpxiP0Oq3efHps6rVPiCK1kMFsuj1YnE+JshAHip+1K3H9AbWxVDCC
meYC+/KTQcrs5+Xfle5mdADCQJqsfM5RPv0Zl9m7B2/1nlvgYhJRX3ZlY55SSDO2nv9sZ9J+DzrV
DhaOacvEyGqR+fUMI9pxsrC1lp9CRKXUrdfExOvCBpve1PvvXNrWrJ6sixg5EWXTFNVPpYTLBSYf
fzAHY9oNzwEF5yNY7hEen//kwu0M7Mom/6LQRKuuZcWa/CITFoSCDVlLCapelnyqclSAzjbTLl5v
Mo6ZJJ7CZ+/Vm60gqMWJazfASLnCPqpPdpunGVXjiJfX+rPG3bgncKhWw21SQ62QVBS+eaKts/xd
SlcM4tGKQVNuh3o/BA9hGEzO2QJMOn2Rdg8yfcT/RTfFcm4JPvnrOfAVHSMl5EyTkfRLp4304IY8
EZpD2EUyCUWBMZ0NPd/ucj2K7UDNqa0MAp4jomHAfUyG506JhLOu6G48gcuvs8OFxTO/8dWyBnhi
tv91d3bsPxluokdYuzkLcsO7pHO9wEGKTRc8/ZX6xRzfqosEDk5nmigpMLu2lcMoErVOmz+nu7Mm
qo64wp4dgpbtWM5q2gL/9LZHhNgALQSMDY9lH5Tu/swfIB/ybDkPUDcrHGPqSJkaye+iL+GDQUZ/
fvMXF6to0tQ0kD1tbJRhPsSHT1bgKizUNmwyhod9IswZ3htMkBjbwEerFt9hc0De4Ww8co+d2giG
3hZWFha6hjI9+f4Nv8vm+e8mlCSXDioLMSkmyqyJJh1RFUkV60PQMUkMpz771kqxM6R5S2eQ2XS3
p+HsgnrNU9ksuyjdw+I6nZufjTgIhqHv9O4jS0+13BPTOX9Akamzc9UkXH7vOxshWLjA46LXPdSU
iMmENwMPb0sJ8b8fi5TAB2jb3qNlUByr0r6Kr1hutVju6VVZn9+yqooEywNTgYSvR7Y/NYGnkpoS
xShJyRdMKWPI6hEchWwWXQsHlokeP3hhihQjnD7OO5RJ1VEWuuTI7XnN+RvwJvQ6a+4jrXr95F2i
bdcqH2ZAk/JqixTvnte4gdr2dh68Lvq7RJFbSH7vhmJHJwKky6+KLBQ4pMX9QaeQg7ljZ5D0b5cQ
g2dsD4RXBOblfPA7uqqnRWZM0KBwtTLFN7rUxH1MTgnA6oKTeJUdYcUQQm2NPaj/tee2xeuvL6zJ
4bLU/LvFPIiroU+JRiI5OUdod8tLNqxcEdaolve8Fpr0pPOAeE2Pu/ZrCGNgHrnpQI7Od2GbrzsY
57eTswraJZ+AKC57unaYt24pAnRuILb8i7YADnl5XePYm9F3UUR+lVPBiUhFr2QUZ1NkweXarDsK
EYy5+rBaaPlh11V83wWFvVWTyrsPnS9qwvtsbxHp8qxbgcjLuyTe0/4Pgp3uQXRWkkcS9fEYp1uC
W5JAmXihZ5r1KMulc4ZyFAB2yA3dX5y6gOwf9RQRA/EJJ8zVjXzcvBl1w2Q19P2K6R2YhN/CjC+0
GAgLRRaxcK+Z5bdUQzD6UvBQRxqfOcm2H9YgR2eBGPVEwzkrpGaVuB4K3eq6sNFZQF/JUfhSkXsu
hAugPI1Q9iREJHFVD8Zbo6LYR1Fl7gjkESvOcVzS/idYJI/yN3vzLmhPdkonIUCfj7T7RX2F/Gfz
jZicygp2mtY/DubzmshijyFI5DO8ybGcA4nKsPl4zAckuqLk9U1OTTPoMxwdhDU/kL0nhT4SYZ9q
fp3u5mgfCX9yz3u4Gdwjldt2fMbG1PbvW5N19HgnipyLVaVNVSl5xCyIDLiGhinG9jZG0raPgaxv
KlDYJpXVbVdREjuATjBCIVm7M4AmjUvNtepBZZkHjkpOYqTT/KxHPQDlAIleMR1LoTGS/9cegVbg
YygG4H1dxVwtL3gimBSEsavsWQP/+rtdIHwNa++jpWTfv2DcTbN9yKZA7QY3yVcW2zN6icCzryw8
KZvDh5RnlTtMviUsxRfcztlHKgF3PY2/ycl9BFluqzJf548pAYBI7F8uAWhziv5zYvP+Q2p2XLo2
6GIeIyCyL222/EV5LUcxUsmdc/KeoXct1bZzmj6yH0Ev+KEQ65lCeqGJzUbnGle86gjTUjOWmEsX
pSrA2F3x+wOtwU8hSYbgMC1NHvmKk4y8v2hc/aKC1PEOSLyBA7oIjJMVRmny/C7KQOQUZmmfpYl+
IeEV03JfWhjO0xJjKUt6lRFySW0h38dIz0Msxe9XBamReSHuacmGxwtPQFGeaQpbRXImPwFUdgUi
sYs0QujHLOW/f1+WlTXfdBsHYuFriMvLBLDIkNbPTYiNFNRwwWAT4gI48ZaVLhqI/RuZVJz8z8VW
ZNsi88SAu3HHVTHZggX37pIbTair5cS/eLQ6U2bMU8SwFMmKZkqkJrXPKPpsuFyMfK2d0ezWC/Bv
aSZobD3N4HDwymbLI2TPYkBU5aoBAKZbaCBo6xwcZqiC3BnIQx6p95aXk08do+o7sXsew2IObtV5
3ECC8KAmYfoZ94r/28Bzx22vb7BoE/s7zXHFxIWSfjD6BvtavmV9tKjWSzZ3aeQzLkbGOb9F4CB8
7j+dCMCUUjn4rL3eHi0MdJv+IFWhiAZYWTEv0Z+zQB+QYHstWxPPzn20OP3eurnR9uAt1FBL01lw
JQEle/s+CzC4d0uiSN9+5L245h9YWIProb5WIeOorumlFhtGVclBScploMMSXlekC92C7J0hX7tg
eWa6PtFiXjCbpZSVjeiREcBDAjAhCUrPV6qwtLgdiJIzNjjIUmvmK8jcLruEX/4bYDV84kvoGzRA
efkyaN+Yed9mxspw3uK0UdLaIyxL+bb0PMXf+Xr9D6PXF5If1oKxnAqirVZe2pSH/u5aQlDmlQLz
QC9GYJIQAHDSjMDUUnbnlkhp63JWqjWu1O8pwkcfpbIK7M1RPDoVCzP7nJEltaaYKrA1JC9r/cbf
JnNMsUjJKLJZNWwXqUwFBYCtBJzLx7OLRt9pBY+LIgg5i0U5kRWLBPGCGxevteFNWWJ7OJs+MLaz
YLd16UY0umleQcYjVHOuymSwI5zfFj1OyPfyG2LQDY44j8jBxiVPBae3ijZkpdLJMScZdbIlhvrk
h9EVV0kgQNIoqjgtZNa0dVB1NTb2QNLZK2k9kG9uEab5eEdM+isTg8lGtvqbwsfr5bG2NOrKa8wV
LhJWSGjAMjESvjSHJX58jiGJcONcWxNOMHxc4C1c0A8ilnCJwo8YUOwbflENzi1eowQse95w7uvK
/qJ9JsIejiWCyCIWSqhUO5+ftUbI8K+ccKUmVmIrvZnNenml71q8l0dSjwVRowpJNmtU/ITTpnJk
4kgPGhoUK2KaiCiUjRqHNeufGgOXAxAjdbeI/75fMJa7nwmL6upWEvFH5SD0Kp2yDYVzH4ewECBZ
gfijQLbeo20GW/wKLOitqf4/CWaFFBdpPTf9UPYva3btdexGUZ/y5Q2Hapsu1l/S9956+NnP2LO3
IMWWWLvSD+7lgckFRHwh8PqHctg3i02g5zAl67LdHitbm9TSShnY1dFdhhUXWunezWuTQFJFmWbA
1+UC3GQEqUNo3/VxXmnV9mfNA9Iq2ChHB2ttfV3EGkzT0JtQpHr5RLPnERzvqmTtvSOYbt8u3XPi
PUsZxMZ+UiScnj7SzyFtjKhOeux/zfin5eNc2vzypTc02XZYs43OK+Kd/n2vVhGTftLAXHQpRuEj
yDmbF8KKiDlRmv7oKCaaO03eLMT/kWCogZRLIuF60u40kbM3ltPVLOBZF79m4rzi47RtSXZ0Y2VR
LofkQEgjj4/EgBvG+jwZkr4EodEUKxSA/q/nvJ49C4L2sePYUccGWrTDrXytlEI7+2NgyDKN8/Cq
HvAN/3PWkNV/EtSHkIF+zhfJVOThRkSo31Y1jCaHnDYZUq7QLi5yME7UtMhxc5xBtMApdUP0hoIf
DRhY5tn+gPNih4ZZ53KM5aIctSmWtNU+3Bs2xfFol8pUmeum5E/5Y7dqqMcbBp61kDzO4AgvQ18p
ySr5ncOyTNNRulN/jmTOsPIRvHQuCCmMzUTVNwoZ7kbywwMeYi6OMsVRnfp3DygWyaPB72p+o9Np
1aF4Skif7lLHW+Dm86odXTmQdCFZyAeVKmi2lNa3ZnW7727EFQ+snnaWyUt1MCYDlrrRbb5ugT3S
uu+QkWDw4OEmEMyalYHamzr+V2+GEipztDt1ZI8utAhrQ/XhsU0y/Jaxypo9Fi/BiHqJbhq54Y1Z
m4DoUZpjO49groIDOE28lwzFTOGQjzo0g33k2Xl4nYi/MgGd7SyvyOgLozX61/DaVBQvG0g87k7b
+3SY6OOVfgy+tUi32MVJPqb6fucythahMKCSPEkGgsE3rrtr419beFbw/JGGxr+GyAP6UhQi9IjS
X0fcMb3QcRZy0Ra/nU8BxyYYX0CHWlYb2cnQ9KpV15stOosLOJbeESNCObjJhH7e7Jhlf9c9rxi5
0oKuqIVnjB9qfz3fuvSVo1kopME+7cdui68uOPLmxg1aRtZJOuoPRCU8IMLos8Tng5KhesKFwem5
D7Xh81xZXKlFle/21CPm/2BITZ+f0kUb0CpZ7NpBu+AmU04UZ0lusKxzHYJ/t0MGcGnCzHyOTNHt
muGWNv2536cwne7hHUZfGoKdB5PRqRd7qhodNBd1qRkf1N+wIAVCQPoLR3GXQNwy5QP+dGcGlgFJ
rY2F6GIspEz5izzPLSsEXBReCQ2aSkKmUS3XexszJieTIaj1Wv+59iPZPLS2qxQ3gbWfgF9WtkyW
J7FC6Bb1vr9a9Fozb40J4lQqJzYcjuSdaO3k0vBIF8RCqoeBkTf7uZVv1NZKBp6M70FBgfCkLji1
o8IG/U9cacMkW6wDEKv0v9o6cH0yTBy6jOGlWDRAWSXFRvt7rpH5kkm4YJ52b2oojzTdwEkU2Eer
dwDS62u+fdXCp/7E7LcXk7aqv1x5ThPnIxoOA4d13C5iVVlXn4VxiAi6kEm1Hn5ypTaDKAHtx5Xp
XbPxlH+sIJLldEd57S1iRFn56s2/JxE/a8tbNB9otsLZETxw8PaeA/SEkhDJXLHMD3fv92l3Z3MZ
U8GyUgXtGnU1O95Na7RfTaELYs/gpCsm1ig559WQIXdSNAwdZISsGwtTHqrEX2IoMvbF7n7cRlTa
mW5dQSCQIcyIErQcgNfx4G6tiHItk0EFmxmv3GHtKI7ioRZPGh9kV3fDOX2Zu2eJUQd9Xgz6eM2B
Dm5DMm+h9uR70nL0IYEoRVwhzBxCAlK9UIXPIjwjdpFcuQRGMK3eAEmQ4QTNULTIKc3CqUqoYTb7
W0/0yrAADM28uelaKJ86shZUTaQjm8SoWd6geXw73103K/I3+laIdmQcNuW0CEPfD/Og0o7L9iAM
ddTPRmKJoSEGcnhJsWNCZ/chQgx5fhwvrOPXmSA5vL90WuzJnyJJzpIfzLr+gd6u7NFhbf+cauF/
zEIX5jb2JL1UIAESowg/uLqzTe1Wl2+JAGkVBKK2op1zoaNgrUl69rVzrtSOpfmmQ8CeILV07aOB
dHb/IjZOV2ukxjaeaMYN313cElXFge2O/2X9YehCymbtRtpzXs1w+JDtbHnUVgmX/XOxM2xnLXjs
C9pbhC8iXmDf5chyWgYOgnLFVWlii+cj6Nc9fh3OBOXMyVWP6DxWmnfxavzmMAp1auf4Ib2Eyv/9
ApW9VK9dfwTVoHm5CQgCaYpOZwOLWmVjoDmveaxZHxlWg8sqwsEPQs2T5C/rAGFv0Zm/XwYOwzjh
SFJFLKhYRrYwRoQgtz/Yf3oTzXGGk6Kpt6W1zhpFAa0x3R7MVHv5w9e6UQcotnIV0b5xp2REh0G8
XK9mBZ0IFfFT/Qw/wWqySowwiLysIIXyZGmB2D2ag7zjLLbjabw8953Jqdjz2RaiAZRiRliL5uZf
l1g1pvrXo1m+Pb67izAPOtTd7FOXRIhePpvf7kIe9T4+rrdggOVRoRnjnuo4MtuTWDB5qb4Aron6
CKP8OJqKdOx12DviFJQdfjiRM5X+e13Zqa/rBKEFhydBrXbCsBNRSRJB7BfdwoZyMreXcJcUPj8v
/7LRFuzdU6K2MozE1q1NxizLvPq2GQX5oWBGlXH1D1cIuObBhK1SsVYj1DXYuVZu2xNRiqrwHtAZ
EC+Mi7toCFc2B0XQ6nO6Ux4IUv5J9Ht4BGOlY6YFhs2Ig64RUOOi/AHbPhcdhsdA7dK7M04uOyTj
GZl3RxWHQzllj5kQiUgk3uMhk6CpjBFIcX06yusB0HFth79GyHL7/Wko/tSgJx+49+fgNMaOo0gp
uXiYYtXIE8memORAltSpHT0qmtKFPjwvn3LpoZtIu5WQUWtmxnmdx/fyebPog8sKY7d9jEWBvjmL
tqrusmJ5RXLCFKLAijPWVURyJIyj2GmQ346J1mcDchYhLVwA2dmjUa4axzbaQN/v/qdtXf72ZPFs
xz2X+l9D4m/g0RwNUffIbbZbLCPk0aJlTQ3Kn5DntC2SbmLBmnfJ1hm7VQJ0k2kNop+vDRuYti5r
Bl1UQWyGoOPFOPue2Gnau5/lKe+WGjnbCF7Se4Fv3zotIdqmFiE/arARa4I0LA+NcNWVwSR5lDot
gCcRdEkDTo3zjFZs3Zhpl8S+QWlBx8iPuIakYEEFOY9x2j60Up/2tjO2FckEbtVxmzZI96XIs8t9
AnVBKgRf+tRePOh1VzCtmgYpnoyk+iW9Y9193tCvGLDuf0pkzXbkBqxAx/9+D8GHHnc8rcHI89VT
pxbbSjOWdD8Mw9d3yURaaWeiLovBmOsP7l30dwK4nscYt4JPDIthP1hgXjdvT973frq2zJFXO64F
9SxfFP1NkIsWtAWhSrelHTMNan3JZ7mSW9bfN7vFjE4t533ZZBsswrRhmObuU6DIRlrhDbvmVxRX
JTFwKJY/mkq+raNDLE75fU54Nj06ezyYDJgW6wwu1zI0dKvZcdRzkD7pb26q4Yr6OehStB7+SDEr
OXw25eRtxm1SAwgg7zVkYm2AA1tABmOzrnpc/dHzaRZ6kxbNqwOg40ScQPWPep01kLSenE4hDAsh
+Wc3QMSSmI9kg9AXXIBfVStRpoEJt78S6v2Wj3U6cNu9f///hMRKyBfYyyb8rS/tPru5pG6AEIUJ
okJqtSg9vhrXPRYclB+REdhnWiLg5AtZgk2ycVxBjyKeLgn5cvHmF9Y/Ye6K7i39XLMWSt1q8s+u
nV5DkdXOMgaVD+2fKjJlBaxrDaNcR8+V4+54dfLPusXYtTugkFzUp7g9kNuQTW+FrvCGJo8Mgolm
dnzCUIKA4Mfs1LsyLuU1/DitHAR2Nsxe5NBIK/JxiRgVJY5wb9wD8boNVRNT/sJXRNVJ5qP0Ixxe
VV6gnSFgarWnU+PbnFr+9uN9r47/96vDBY+ENrOkpkLgFmEEaUs2JJJgUe5kbb+ufh7OPMnkgoay
2hdy2TOKRJSbZtiOhyvifNNB3O7Z8Hy3u+Masd2yy2OQ9R7mgC9zBsrMJGz1m4CV6UoLOqmBuc+l
gaKllPHtYbxF+2/GGCksnpD2tnC2SgxHMVqkN8OedZS84KiyJp6v/lDN9Ma9oJXXouUhLgKQTLcR
P00iPNhI2kMfqnF2oHMAyBgdlYtXIpOqwkMmpE1SlS5aOt7y9RPvTeS7AoTiItuVuTXQ1obdXkPb
jHfA4vFWmsxpgoevCxM+YQPNmdITjmfP4saY1Lswl2DOwY+yyAYqsBYqxXGhWz0fIGkOTFHWBuRY
GezYC2zMwillvyMZi+j/HOU/4xOTfh91dT5sWrbyzZaHoc3k6GzKBZRQJ4oFT+i0kxjYilXngQX6
xSpc+oKMgN2fyxPapQUevwgpJDQvR/BJAIMsd0umOoiWgGhbAB+5aY50r5tXWbvbEI5XHCoQGUQW
ydh2tmxZBSXl3vh+QDC7+zv/YoXnEbfF7a0ob/2vDQMgGayVWliE+knJcHS1XBEkSA6fzK1sYQcj
zYtyArpDiEJwAV/Cri6wCQNDhAN+QOSwIT5LBJmos10UnrB55/M21EoPtXp7b2B2QF5i3RizIOlj
Wpu7EXn3HYa4BLptpxw+LrrX1ZAp+hS5vRubc8OiihlrDLji37NoLGAgKEgFxhiDmS1FK0sVsFBg
dbHWd0WvV1Ayk4xhLdpA+Wohn0javshJ/49hgegqvy+BeZz4+eTkTNzi3qIjmzDjbiUTDIcVyqYJ
KRH6I68FMwSI7czBqhsB9rsGusZFbAox2xbIn+0bSDC1mJCOVt7Blt5RL1kfSg4Qs1RRiyElfxlX
FBcTpG5/fYW330yFsSB4wsM69635OXh0RxLxxcf9iMeWhH7hs6p4L3UX9URfXsOkn/klLzPc3aoS
HrvDBmzBlYkqWmwPF9fyI8yVa8w3OR8PY+3IewVNDp4ok7VAgY3kUYeqXyzEZQhXhB3o6owwTkUP
F80tVTlsaUXtF6kRy1pLvBBAoM1LyvCNf22627sIlcHtRoAFlTmwEgRJ7vu/bcbxj4FCtURwXb7K
1UIpxMex3Q4ktNDU73DeLTXpiyBhEBQ641GH2PabohmEgzgfcrmidZrY58sM+UDV1OvpqHOaG8MR
J+oJPUcnvH+xJSeLoBV+JUl4g5SYPqS1VcyV35Mfi2Fo+/bvrBinDhRP+gx9lMlqy29bGnrziIs5
+bfz6mxc/nwD6oAlOBngYtOfNzvy2NVDAJl5jyQgnlbWh1qpAKreJdAGGlDRhBaANevEa7D2s1sV
gEha9SGX7f2beNFrUf5RW6EJSA65ue0XjxlhcvupbRO4Qt5in5XSRQhLzc5S73F1V5JUlvoCojpf
Ik/TFZEOXGLN8Jc/CsS1Z+qF2nGeWof/u0ZbZDASOtpF/pvfz1RcVsX2ILAdz0GUZBhj12MlpSbt
BV6zWKrnIs4iP675dyd0pUqEt3lNb1ZZp7athvGezN0dHeP9PQ+XNByJw7RiBqnDAjB5/sNVsrfn
OTYDuz7QIdmHfTtsAmNdKFfSM4i3dyyUB1gveefKoLtisAWTpTL4jAKo/+aQc3q3RrY8kUe8dAb0
wWsuahx/KXyIJfpslFjirHcd7KQEQamxZ56txuisbgE9Wdsyty8O/Q+FVeoqCfxpCMgtxTx9Lxjx
stfHB4eFmGzpALDUGs4qkkkEGtIhDw4UZyN2ctv9/y/Txam06mgakShWElKV8dyRWfx5NaNd6ZOQ
/0K4nDTwxKOAvv7CK7azdxiC8RgmVhMa+n/anjtLy+0nBwahAiwae9KExpB9vCEBIuLPanjBr1WV
Y8fya79NiwDnXbflAVqfJmCsKnu+zC7lc8pjTjZPQqDSYsnaeLaeOMeZYvnxQ8V3BL5opHUSP8O/
k0LB7Dna/LN5PqI54I5TAEZagP+BVbFP060CjRF9tcxzUcZMz2QCbogRQUDQv4Fu+MMEoLABMDAY
JMoGldNLkE37WJN3/AzlPc53yEbRa6FrjRCzaoiRPrsLWzzVYW989YO9gHHAL4A5VOYA20OAEFhf
J3Ad9Kgll+QXUEKQ/pqyulj+TrIORnXeG17Q9HrlOQs+Kr+7QEhVHti5xMJ6jaRO8hSyDFuj+Fdw
l9TeRIaaaeSR/eFIPD3v62H14wWIS3Ky9vqY8aR0gS36IEdxqPtvOAAqapZcPkepAO34w3XfperC
tBgV3VjyvCB0AgZ/06OGpE+lDtA/b+MRrcGEh6B3fc1GqKGtyRvzH8Y1e2uJQs0guc0x/WX4R9Do
yK3uircA/yZGOGz4trty0p40JF2vD/Hp1FfzzuVRApLQ0eizHOo66tgAjkVos5BAQSvyOp6FUtQw
ijMbDZSq9k57hPT32N50mfEp5VZHqCM4QPn7fMU69k9oc50XCrT5vzRG3uBu4mVXg21tWqduxY4C
W1odcIpmLBjyZuqsSR4j7pRP20J7a3XHYs96tKRptTWVCal63jWcugE8tzjI4NTAEqJViViD6dlL
+/1g5Gfa+8/CGh1F0ayscfvUaY3PLPhlIv4UeM1BZx8jto8LuI9vWgkYnS3oCt4bk59AcFNptLBI
sB9uFEO3HPdJATFjAuBri7BhdB9t21z2yqlz4/QttiaMOTw0MlLJ3nRiiKKebzfrxe5FICUSNPBL
IgE4aMDwqbsn3jWAvSiQImsmbXOOPz3Po9PaABEBb0MXl1oYfLZ7HxeDWfb8+EHM8dvEPOBf2QaM
o0PKEcbYbw/pSQdZm++DruGC+RZliKhH4JtQKPUig515bI9pP7oDMDqWqvri4ZQGq2e8/r7gjyfM
5us76seWnENixk8f/m11WFn7msbPkzJE6htR1m/eLvuJh1bOkiaumMVOEIaz4TsPpB6oG+DfeNeD
VUmg5nArCG4OAUfUCmk+GwaoNni3KmwlEAi9gsf+mKfNuuvwjfX4Bnqdz5ehZOy5XQZjONMvp4YZ
p64Dxg7OxW7fmXMznQYI2OzcMHVRS2pIpolPMFov901MeSQXCq9hbC9RJoZq/FN3jVVLoM3yvb0v
kuHeKN0fdy2OOKDSO2TVumCbRpwDY6u5lcwyHHVJDpRUevszG4QGVPxWaxcvVbr8ldWvEMW1eAOu
qB5lY7O/ixjcBt+T4mGYIk7EkBa8aYJxXynBnDYGXxyGCD8zPiQMYqwpv4JywwSGPL32dbBWDoZ8
1eW9+WHRsbT7uCV2Th8si48K2bT4RWN3eHQ3qQQE8X+6PtOkfwr3GE6XACludznMf44tuTTiTigI
Syzk8WuATbbenbFEUKz2QE2AojY4zDGMA/vfbus8WGF19FViodOmo4KxqsNwVd/20Cy+f52wryhD
XviQMVfuoiufRvTFCRCdkghGvaBoo76Vr5kBCoH6ctdzdWSlrjRzom6mfeQlnaScW113L6/dTzXC
hIBywl4did7wmjFUIagc7PoY+bEtj/J/uAnMRaND1BG0ZJUJ/DLVcAahfjuyVu1UMnIOj/MdHEt9
lFASEbsGCU9lmcCDzu9QvrTPxYKksTkm5b4KE7s4th9f3nwg+TlBS0gQUmea3YBcTGZuxHx9c5IR
rZFS1hcMQWgIWERRKoQZFPKgwymSBBOlY82OPzPAk1bA80Yk0YwAknklEZXFTrvtQXSS+1O6dJX/
C/pDKunvD2oMJ4FJ84OlSbMhRwrNDcEXVapCCqftzoDKcPinI94edsQ7UNjnqRSFrVSv9yJW+cga
mvuCfcCSVjSXKZDsS5wkr4jwPQ0OoeGjLNCpe0/uNTO5TqGXTvo6VPQ8u7GJuxQ+5L2D33EL6KIn
cDNjrpCPdz+3E7NhtfJ+TruYztubodNvGvBAaFNxWAC2P88BlkVCdbRSgQi3wbWW05HLtrcAik7s
gl4kymAjO26Hf8mBo1mNa/xaBGCT/brZdmjh8Qjw0lF4OS/h4BFo+CsPs6QANd5sVLOQIYRr1+ne
e+SxPPrMNlKWAnFZgCONdmBFuDQ8j6X3QM93rM1dijDfplYQ94HRDm01QN+q4NRkjonleGvshw7F
puTDv6eSwB+sWQuntwj8vFmFAEsZNRYIzzA6kIeVtHJnfISyaHhyEb5uxmCMmt3ugWyA8yMB2Miw
1EQQDgScgezhWtNTvIOCCU1OO2zYpmYo7DsgxvNDZnSupfbg37g09pAG5JnYHaWvnFgF+pJOU7/P
vyaziG/mGJjqNMNd/Xv0EticUDjw78EmVqpbVcPDUPT7iYlqaizVuV2fqRfg4pXu9Zh7RkRyP9h8
vmVyKRPYv8L7qmSkVMS3kHaKUTjPdWrlFMj8y/LrWqMwkmbTvMHb69hlCeL+Q3MvC1p3bMrCJjLH
Vg1Bv3A4i9iRTEtp32FFYQ9g7G1W1jnTubLh1Ql5hwr7XZeDlrdLjlWVNxwxovoyLzHGbZXshvxX
foHvetgt/UjgwPx/Tt1Ar3TeIBLxE7xgmgpfWwbNrk/pbkrDutOO7NPpMA4QFulTxeuWsIs8CPVx
XrdeDJZR4uzrkLZqONYzpeIXu7Ka+lXPqWlg0rz97RzTXgyonaV4JGRpo/oY1tktgDnZ72mT+Py7
NVeuPM168cLy3bWwlyaCqWKI8KbHr4XCoSqwI7mcd2LsZmAzdJGr0eVrnyNasPD7qO6+V+woRunx
S0Sg1jW7LwyTcJY1azQuhwI67Bmh7EI0/28HCeleJbzRi6+aiRw+NgydL6SSwRrxF7KzqRY9pDE/
FcVvq/ztd42e0A7FOidNWwUJg0r2AyyZ/xo5yQal/bURzNf97amBW7IT2ClyCVA3zAIu/zalhB4w
1yJxXZtzmt6hiEtMIzEFv0mz/RNy7/myMue0Yf9pIO8Ia/4HxIpAwnDs7dbZFS2iyvqxy/QpRCQK
zTDnvqSIF6XzZPzVvVp3FEeUkZcANjxpbuk2qXk2Q40WJFKEkWuhrNVHV+rjl4IeNfuPhRmPRtDz
rkKZFTLepSM4hCw7fo7AMQJLzN5sOfGGL9k43KXM4aruTHG8Stnx7yxyiR0BgvpZoxJyFV6Lzhhi
Aib5jCcwPaIY/TGdm/AtoJNFFatx9b6Ln3fmW5U5VqSc5QcaxXp+8RstxR9zmFIW8AAo8MOi5XzU
XdWeGVaeC2P+rSsRjfelTog3vn3xhbb/l3aT3sdr2SHsBb+KxBuLu3PN/Qh4TshzS1QmT5UmXHBW
45cfrtjgX4BQYnH9jXwOfxaqAOWbJt9Cym76LqyWEtLvy+yzKmrQAqPqSayS9MxCYzypyccWg//5
3df5+9d+XZ/vnnQ5FzAAQI3s1cY0uTqqCwqqQOMC/MLbuh+/n08DLl/qFda0fBm5XQ2CT5MSw3jg
nM8uM+WU6Z/9ZUSJhdHbbvivyY4erpTHe3brtwGcLx0mTxwNxzFJI5zzZnktTAtFelhnmqWj5FRS
XsCb+KUFdbMDCMh+bVACik6H+TOpwBvQqPgGEvDL6+ojajk+FOoeo2xxL0CecwrQrWIOyhG52qaY
po/ysr1evj/C4GCgqDchF7xaPHgwuyZz+/UAYfe18BEf2bhfvvpo16ROIx2ChfFV6sVNSUBVpbce
6h2eM1salrJKJVXkMw0GU9hskaqC14TC6JI8AIR3B8iAY8S3v7e1uOxOpRT4l46eU0B4mx7m3y4b
zXzNnNTSHfh9J+Mp647uRl3w2RWPnUFGrmpUMUFoX2z+FvzAauI2wIdayvvRc3W4wSz3ulEMhjWa
y3Z7HWCIH6WY32gNhSuB2h95UzVvdMg3lKzk6pWCXUZFQCuzkZ9MKJFEPSl+YgbTUjCug7mj+pRt
3p/n71ulYM1l5dTaFLXMxFxW1Ay4YQT4aXxBDl0Kk/39gUvaL479frqu1Jduss3cTPUJwrMTcUOR
Fgi7f5+VSlzUfQlW4pvS3FN/aGrK4BnyOIDN7JAjz8ELT+ixmTv+oBCqkS6WvxgjV8MoNrkfdMhh
e7/lIqchA/vcYsd1sT/taq6lSBEB3HUc1T6FoO9C2xAeERiMt+c1qDX/NNlyBZ+zBYcn0CPujCA1
OysZUwwPk84GQw0w6dd3t/ZFAaxgzTPE1CI43nPXBoKtX+gABNlCqCp2d9EE07AdBaPAx/rqA1DF
tIXl9Wo3bW1MCJ3VfENre7seTe8QAPH15i1LeAM1ZaKj+yzhOoTSbzWAgxJvzBLdcfnOBiW+grYr
Xa75Ot4M74VcBcoYOXLT+vzvIqCvTBcQS+OWg6vqHiL8SeC05+TPrPAvRkXFjVOH4YgfwNB4na09
pFwgCcfLObKi65jzXQx39jA9iF8EuiR95wWWK+v6abnjB9f/k3A+nvGYOKuueun0YSrTE0HPaApa
cJToFy2VgZ6dvAdkI2eeXNd0Uk0cq7PT47vO8aDplM0gXMKZqKRTFBBazQlCTpfh8iFHgqg3baTd
dmk+J659vPMZu7BHmZKEmPwPV2xBxP/Mk3GFXKOzFoIdlCbszkGU1Wdw8mKZxC7ngPgYx+1kUi06
k03Vw/MDy8dKaluzx/Qrr6crzgoXObkk3awf2ENywvxo7SwuNzsaqJzmHixt1/pzw8GNo+gbEjdR
2pC3yM4P29eHUVmW1aMl7G4wLRK4sSrlSqt8ofgBmuJPxZIMDc91YIOvifqQ7OaSq0XEMJlrXGiL
a5xWZxGt2v8Mij0A1vFlrCuAizg7EiXtiXajkr4nlbaxwHa/uY6xBtzXGkvFzxIRMC896eerWJBw
Avv72Vw/XZhDhn4687iXsmVcSsHCx5lo3kcKB24Pi7b+snYtVQIt0i56BRiNnP0hlvaAVJxrJTvj
LJxHvy7UQQDObDSpPKE0IM/rgm7J9X9oGhgAcKXlazTMZHWC8cUwmrQ0iHAmot3xt5gR3uVtAXJU
4ItfsLLnI6AmdBkAGGm+ihPTuJITY+V+X3kUEoxYictIJSsT1hy9yC2zl1UQJHSQxYKR6AkrQ9FZ
Yz+ehxASTB9YiCtn0oqo7+CtAOWOFCjINj0l4CLimxU3m0RRXq4d6aVW7uP4pzlHGa1v1e+ugxrZ
c8AFyOJpPDV45W0wDfN8ADDQX51wmtdpIVRqN+eHx4E1y8XnTeWkIGMfXukrREmBNt6x0de0vAye
7cJloXZeu1dzOLgVPZyw3D2Yz8CPCIwFNNhkC6l4JZfwq68+4CzsOQQisZipyPLq/qM6jJeDXRF0
WrLjzt21CKcYj/nTmqrsdFJOEJpTV4L6dcF5XUVbtraZexJxVYePFNCwRkns1r3nIq4LH5Lq7HPt
SURjuPUGh7eY/0CKaMpSh4/lI1OCB7PDrGmUtZD/ssTadDaz8SCtxoOxrfCOP9D3m6vOqftMjIae
nRDETejAiHgNwgcSE583M674c1N11yJhiiPiviw7K8QlYTo04P7XhTaN3En2AZLOuusuUyd/iCRB
Q1Orhmc2eSZa3xtLoE4QX9FcwNfqlqfKhljXs58yYm7STX3Plb57wWi3u4g/I0giCmK3S97WkrKQ
hsOB2JXiySUU9qknQfV4Fynq23qj9sQW2mJV56zMpxK0OphWEZesVv0NEBN7JI0hb/C5W7VL4cU9
kCVFqqeXSZjYjLcL96D9YjcWJHlhovVy8Ff3f8t6f5O+BemLdjPgkXkJWUytOb3lgKcJoWLrJv/W
wlObSYyfENBdFYz55ZmnE424UhR7Uz9jVKL/BOOp0UkYs/ubgBiMgcJZJWruJV9PFQKlndMB2K4j
xrMMl9q83T9QB6jwd4cyzAJ561wzTSkrYXEvGv1O3aXQL+BBSsv+eCD1xwviza6uCrqD+41ef14Y
bJ1+WC6+DOB91uiXUi7nkusuo+rHwdiZJzzqZVYYdN/zmE+Vee61b5LuDXTzXkc/BQk8j5oEZyww
i8Zh5dlRMLfyIpIBatK1864x9QC68EwLe2E5YD93nhAY1VNSQa8us0UuCm3lMQjCvmdYDh2vGpN1
+t6a86XppljXLqVWNJUpbtl/vj4z12+lW2N3VbkuhlJb39KNZIEIJJUBjiOgGHRMYJzcscFkfYQ5
e2RcIPAIb/XCB9aY3WCIQhcuSJ1SCy5Z6TUPQqc9T8Tb/L3Bsm0tez99SVuItxdnqQ6wnZeeqObT
P1nNthQPKpF5506JdFt3XnqaXe8RkJRk8cevXtlS2vJMjCjD96ch2zoeAySI8Un4NBFUQEOb4QhL
91IpNDdYUr8W7UvETJ/7AbNv8BQVFG/H15MD0ii0MWrHvZaJ2Nz1DzxzHP+CTuc28YMUaJ2ZcU7g
0TVZ34DjEteF9v5hAwQFSO/QlrbC6GVGPXwgO9RbmDfL4p2QvIYSHuTp12e+m2VNcQ8zYVkZ6yb1
tbBsH/YMqWWAUnY/iKiUjHWan8WWEpXevVnQl2FIusfmj1r0BpcC5t2nK5I88QLvoKwQEbdoio64
6RhFkmnI8EbJdUEid1O3HfqMQDwleiANshGkgBi1tMpfpwEAk1G+XFsBtc6QDkWfbaOALliaU55I
K1IEcPJzbE+WT5sDFWTV7HvaSEotarKzd5GiaKhmQeA8JbeKJCGpvoXeFr60b03YQh0dR8u03brd
HdC5eYGUx6iiC4oQaw4as53WsczE+eT/XlZktQNAvq4g1KwPydaYjG0MOVpajRKmhWIsZrQS6DUK
gOSIHmsBdVekkUJkGrSXV04yeGmsjWc0TNWTV3fMBMSk7OXraKxcs6ssjH23QuGMhwdhFuPcfihl
4ekahZnaESE2jF/0kP6yvegJCy13MmTCLqBhNFI2CRmHbd+0j6IKExOhuTiWIz3gcd18nY7o7BEX
uT88qR3t+iaofVhAq8Jq+eHlLLHxEPe37Ddy7UXFWMcNF7hWhUDWUxC2z+eY9qHX88Yww2auO26o
+/O/4n9AN3C0UImhNhtI8mnuWHEzhmFB9tRm3wKRwDoYSKaYgWYV9eFuWdIZlbKQP9KWTd1Vbfnw
kasfNYnzWog1vrW2gNAHh35AvlJDLqY1J8hS6qTJJjehCgUwJO6S4QI8Z5gwRWl5Rw6G4Gy9hBgM
GomydxrCMydGaKhcz1vc+nEsvoSXiNceV/L7LQlR7NlpjU5c9B+TMdnwrButvAqYdZlQ4EfmaxDf
VxBA8RkFQ04ABE6BsjVygRtnB/lEqhBWwlBJM5lg1DK9lzBsiK4FGS+b+eTWMKF8TV61vFdeKYgV
L1QVWThn+HCa7bn+/LJX4qO9rUKdY1yXCn3QCC5UNMv/NXL2l1DUJoLOXXb73gxM+K2Z6Y2YxRLn
rCmlOoytCEUAJCb9K2s4RQAEjF7KmivVyiVXQjyWpnWir/m586HuLvjtxEAhrEBzlS1ZTqxCxLXH
P2wGp/r1e9cHS3Oja3Y9G9UHfp3R4KxUJKaMmlvM7YVUGMogosTaVcB7EAU28wDnGlm5SjdB1G4X
WD8oeSeua/Y1Wo+tema3cwhiqNMyNkpMAx5YrljTkY6mD9jUo0KGzJYDQ3tl8KOvRma07OF0hn2g
x/rCgN5nliaC1iHpRS12jxKI12A6hv/trrcvzeY4FQCOLapuUhcbeQNG+0KyYcjbxu9BxqKeGHoH
aPd4ZSea/y0R6Hnj3NTSJd8RRjUJkLcjiyQrqJ9izGKABYdncVl6+mSphMu76pawpXRuG13YM8o5
EIjjtBdgCwLlJlLyG1Necx65z6SmgYWBCaZ0Ax8SxmhBEYSd6Q0UV/1mZuQtvgVCPc+awpmyX7/1
24oL9Wg0k3kv6rJYlewsejanwo4cd1g5l54q21f4vS0haokaH1zbA61ClrIbrcUhhnp7UCdU5TII
AHnQWdlK0eOulIw/y4OiJ8EXvjLpSXdDiRPI6oZbKifujTKrzbNv3E++nZuE+1kQEV0ksRw53o58
zs97d3xXOfRaBYPy9Axr3chm4+OeNFxIPabfmSGSdPrivum2/bIC6uKadiBsBf6dGKpS/aTKWc7U
c2pMhgIxapBWAnWsU3v0ps60rCYIspbtmUiL3zV6iB/5WHmabksSAgzG1BTkV2I1/jxohg3NeTJq
JtUaLkqI6oz7HPWRiZl6Xy3pW/n0w/g1bhelzaHgParMHAK6DtGeKqtw5a+hDolsEOicsipQFllG
tw3VMN1aJI+H8J4vi/4J5L/UlgcA5zd8f0P79LPZb3suIPkvaoFIvP50X+whM4odrp2xgeIh/5Lz
6R31cohk8knX3N+PXftPA8XgML0tMah/ZQWU78JPh5AIDc44BseHwZBNF3+RRexjj2rQRvP5h/rj
aEEtYQPbhMLc2dPkdovXF5pbFdF/K+eQwfP514K2UxVfD4Q4C/bNq/PAtkU2hqsy6waTygRio9Bk
UmpNM2kbz+aRt+8H/v4Tuxtp2GmTj0qspq4rPHQyVsgnFRiBdWIbObEPO29Dl4/aHYA9OW7X/DbE
UKaQQ1rZgyd+rSjMQVa82mqWbXHtLoOCzc8jzMY2V1OwL8qD303lf20C03C7Yy6vjdbdy9u1T46x
9Ebo3xLmsMFNnZeZCw/odf/z5x5TzymaDEE4g4a+uW7Om/ITPEjgFUugcw1sNC+Lzm174kdI6tib
5609JXDDpvFqaKnwPKPSaYL9knNt+8t0ZAl2QcO0O67ACCWS4OUK7WTcBkRLQhNiss2c9xQWAxPi
UsV4a1/pkZATgMCdYE76LMt4pbvks8i1C9n3xd7Gnu9US0/MvfaaPhuDTuYB9gqs3aPPrG9eN5tl
3jxSOr1qOqBuTnFuqdYnJquTO5NIywGK7doy7dGZGsZbyLsv7z2MJO43+W+n2QkcTPPyDVPSaCnE
bWoTC6g3X7TzSup4LpVgKZLKw+7gten2WGAfj6zNl+W9UcOksiVV4Bj49ENpfmhOrZcp1JMQfKDn
Ymxc8jvNVNslrRlGQTwtSNi7Fr0DPRS/tVNz+l/ovDSkLFq+AtVFolQ6zj3dQrKsDBhe99nkIOdi
noFIFxtn+XceAhYgiq8oWcwkAHu/N5/2uYGEjOcSb9DKBZ28jatQAaizkVUUTMybrYGvgZKCe4qA
EKCl8X2ccvX9zlP8Y0ciujAU10SXDz8R8vssWksYhBKqRawI+Bon3nDbM/ifMexhB3Fi8RZpFd7P
BL1Xh1udiCGwNXazFO/WyoBMJMIfJ8VzOpQl0FxDTE36IWPHcRXaRWVTIFIYg1pbQ7fw6BNOgiZd
iKhp37hD43zxyLMYpsEiprQlvG19GXGowjd7jENyWnDXFbDtkYnprgttxLIei1nRaZVV+hAaKUSE
HZEDYd/0baouHlrosFMyxewWT9G3Mq8D2kukrhKGY18s8UUW63Ol9PLtJ9P2nNqjIBAYXsEJkfhf
lrpa5UYPXLfJ11F05ShdEaCWbgnTflww1C3YzQJX8cW9z8XK5gbNSlYWoigj8eV7c42LoCNl/4Ua
mP1M/t+u9zY3Sdt5iFRAR4dB+xP219yIApuzbUsq8X5Z3jvfy+/w6Vw7PD7jINFC3ixvSQ7q1W/c
jjOzZ1iO5mQqIzUzVVi+ZYWOVHXjeCyeCGeTPk9bWYkt/ZMvVBfIvMkRrfbieaVcuhajT1VvoowQ
C9pgyJfa6G63bfU9Ja75sie5bvSyE2b4RryHYGZMhqhPeWh6jFlBfYqaPm9AQiGlLVWS6JOdqWNZ
FvaWAF7JHI2sFHPQj58DInWBQcyGYLHER/b2l2935tqZ7tMoaxU4zR9zZcULYjUGUT8QScPdaV28
Z+B8FGgV7xHml11tQ4Sq6+YiYbwLegUicGLz+gtnGy/XCYCEupuUxglIf6UOVAvIL76mSHRQsg84
QtChl0TEevJyzWCmi9BBJcu/0iVqkPkBUwSk2g8U/XG39sJN2ZZe5JjwrrTX1ha0BFjzQC58+xet
yxvMUxpZg+NNYuJQCahSV6EbMD7LrhZphWI27d6aMPFZ8AqRGkcL6CjWKS5bx7I138UnWrLieM2+
bJ6XiyWjgm0A4z/4LOf2DFL19rtRm53NK/rrpAdPk7C33lLeUqbjSdzksiqlP4iAkWYe2NaTkYme
XvTItCEw0Q01ANAa0zsWcdkz9tYbjLBAfhB9iWjVNLI1Kl7Jc23hJL+62DwtXK2giuhjq7BNfFx8
/FOIvx3p2UCsOjv4kELKxgvk5EPuLeDYiyZJ00jYCxCaumG9PmOZ0BgamiAfDqQFThSWFjmOhHNo
WVUJ682XKlf+4tg0UudcUqHdb8UFmEtSgxdGtStzcwe5uGXTDEd2IilYNBVCrslfUBfnoDV0W26n
bjuiq7XrEk6f/iHU0GMOXOZ9y3SpiFJdCSg3BDI8rNi8GLUO134OM7NEt79hI27CIws3ne/cy2hi
eGjXSjyiOedTkg4NZlsIbkxI6IJsqI1LOhMIk0mm8tjtVFlUEb16wgFn8LrJcyVEeUgSZwaHDEQx
HP3FPl8niOeQqL2z6NXAirj5U+14F5MzigeG1Ja2csmANvipL75sac+evcd3p3l1b/pyYYoMVfNK
th+d0hcTMK/VnvJAGLOgcm7YvmiPcQHWZxefbVTo/43cSurzXFh1MkWxIVAV7a/onko0IMdqI5+q
o6/6dszhUoCf0U4e9MCLx77EQtjerxnwBE2dkthjCqsQp3ztoil/dtmUoMZCe5LUcIsy5dIi7NWp
JemjaEobmKokl+PqD16Ml9yU74YnaPHcuD3+07phoWOckF0CouymCZh9GY+wKGHfqP3nHz9fEpBK
KOersYf7uZaaQGhxAUTA+3dlJGjHhFAtEmmq/7bsUMPwsHy0MJdrwUBsQCVPfaQfm6St8S7BKoXd
Aib2Mk81kk95qn3BskAydQcRU8NtWQKjNjHJrd9A62/IM1Pzi9NZlinkw3uXhQ3+u1aViVzISaYM
EgJ6GAMkTjx6h9G0owgFc448Dqi3EmG7MoBQVVEek1mOOjxv+f4VF8bvwa1+Y9nUyPwSKxDvtKdT
NyoVQjlsgdYBrWCjg3L4KR7xLk3Wd8zYwsgph5VvCzZlthC99KuDB4m+WHJG70KdTvFHCCQlAF6W
aScigWR6T0D312el3zs3xA9faOh6Q9j7BnwHPnzyZV8tq4SZt6N1bRuYePwIbKvjErYly8APjn9R
eVW2Y3R6xAQ2Rv1q+qCnDxTbFrg/m6DwIMUhJ8TAy+1RudDv93KS4+unOrHz/Yi46Ooe2AOi+vdw
dX1Nu2dEeHVjfObWDkMyQGNKag51YRlEqA5PXPB0eSWTos8OZ0sQwpY+SHjOZGRWEgHOagn4Szsk
UdYkEZxllzmVkPDNzbITPD4kIbcxN69HdSPMWmtJ3zohBVF2aMZ0rJd/EQVC8qySiZsTQF0fkitE
8xw8PnJYRpORiVyWNrnyqqmDc5gb0PufR97qi/trsxfoHbewWEGdYXpqSignjqAPBx9Lw2CjFBZP
sHYPavtjWr+I5izD6IcdAHHjBYKXFkyNW+MfAU6vCvT1ls7zUQ1IfpEHJb+iveZIFJjEP/b97AX0
R726v+OLMIvV6mIm20m+jGJ71qwy/7mbnFGAG1he8JVTEbLbdeCytW571KLocKGwCK+PtuZY3CRt
UmMTVrc5yp7XLZyrR0+omkUlrFT4R6X8DxSovbULDFxGGAykN1+o2sy5ki/0t4FlOiszknnQ4yRh
tkq6K8RcnrgAv4ddYpAzGraTtGNkMbD85AkAsCKw/EXhqYU3Ng99qlotOYFHQYdttV/XujuGUcaz
LsPqRnodRD0+R2mtGBqXzlShaa9Oduv19OR5AlVR5pR8r0ILjtotx7r7IjuxFvpG+8jdkT0PqJ+8
fzc856wb2WtNGRd41szOHW79UbXRJSb0+hkIkcMPB7a0ny7qqhb2jwIc/u3nLVhyvAZzFPP4vTQk
gt6J/zubkJB3D3Q0yeEwAKeAMQdftQd3KONRHcIiQhq6Z7tRJ66IWxMxF1ILG+IVRnM2Foe55XS2
GcEMePDLC+n5yMlVUzuuxPakky3R9RZIdSo2TMe9xcTuXz0ukvcvmufyxBQIk8Ay2FnFBC2rUX7J
E/MuwrMRNiSCoz0mxqlAkZ8dXeLJ/EjhlP85E7VRH5MC9Sb15yolON+k3ECKmqfm5b3VnV8XxQH4
BrkBG067rLunt8KoxRcBvRhmleVQ4XINUFJoclPAklASDsfhSxImDs2uVjVgEm3hU4vlHOnskZi4
YqwDzukhD3GZkzRgu+AfKN7nBMm/gbVlIiuIuPpBS3LI1PPKDp52iv34pGyVMLbX+fpQn52velqg
l8H21KHKX9hJkhWDx6x5nYMDSevijPojJ7e7zQ3pq4upioojYsuQi2z1ie87asB96wnygG3gWxmB
+taiDCtKKAOGV8DOua67P27+rVA8w4CJCOfFqVoPCL8bd8+aEDCa3XAis3v2gSnBDnVLfWsVzPfq
xS1cSuiCkLuTl3f3KBV/IN/i4a6o8MIAzCltOnHS1IWMwRMGyVUbas4rBUGcU3GycnbmsrPKaiNT
08HcM52u7TnY/tSr8T8ie47IzHY4yUL7TuPeEXslMIBbLzq+5/veTloczUq2E2L7bN2ugQvP7BAs
O/TSXeN1LuycDax2yP0OG0jJLzHrAFXjF/E5CmNYZuEj2qKxIW0xwtoayk2z9UD53P6cBydDaluD
j43XQkN0dEZyM9xpenOqdXyWeuqElxR09lYyvbYnu78iB609t2GDRX/OfgV/kYcH+OJ0vzI1+ftH
h5+K77vSR0nk7ibfCX5NBxT+iw6eYWaqryUCoJIswTu6B4VVQ7iMbOoC9YviQtItpGNgvFU4wUC1
v7+SZlU3IiRlXeAV++Yy7uGHAJaiXFVrd5Yd+GGFX2DrHcSJsCpTI/RVYrTyl3vuECSlAyq878Ys
+7dy2I0u2NUD4z8JRdwBjswkY4eeLTo+Oyy8hloSdmQ37D9HG34ohlOLJRp3HMTBLziClWzGgVJv
FbDxZdbH/3Oj4VHvFsxA1J8t8crV1wTWG6pNzTAvWadAUfHWlPs4PgR6ZvXJPVJEM9dL0aU6zMzA
F7JhiLPavkONQvqlBFxzvzlMh6HdDPlwxobBzbSzdd5uXFM9c/VNtIZ7ge14UsdyRcS1xYdlYsgf
iV44M4ql/ayRs1sYE3AlltuaeeZdlIxW2AvQVmkyWSJVQhobl+wpE7W535Hgq7BjHatZdrOfweNS
1xmcBPn6X4kyWgpIGLaLX50SOUSAh5mnYeUWbIHu0GuhTOESfB98CFd19GaToRll+EP6LG8RHiAn
BqJmKIHNZiilCPEOFE5OgODA4SG9E03PaPE5m5GpaiLbNaJPhgOygep5jMM37c81zfXooGi94osj
gYDFzZHgPYY6xNNJx5IPHrHZODp4XgzCpT8hygWlkojhF6k7o0H6sKjwH9+5PMr4baFB+HofvkcC
5gxRaJS0YAYx1whF0qeYVSHKE3L1t7tUMbl7L+DqW3rG6KvjdYWKsuP5v7b39CMeQGUW5FSVJfcy
bsAZ5SN817YboL969L1KDRgnqzFXeFjFDugSLvSJzeE8hk1rw/JctXnqovwYIDmzGw1kiFd3RK/X
dUTAb4hQSdNf0NdVoiKxm//LA4Dzso3mSXkW+nr3zzbIwZesNNkTc/HATnA/vRXDxWy9F0XjItD0
LwfGQdK1qDzOyC9bqlxSAsB69nNkRoUvJctyfH8e6MEjYZV2shq/gRCPuF1F3WOQ4ILoAYYn21Hf
SNgvmtkKhBWo+IHl6lvgkJdJBD7jxNoIov2wdcDkQwjRqrcxt8FPitZHMvBPgWiBToC+szqtC/fT
YPRy2zL4TYHlG5gD9HktUiIoxbl9k92wPvDM8eTNBZp3RJyCcUmbOubeap1kV3kvWj4w+yYKILO1
ZNapXHkXEhY8Y+2DW05LqXWjxCCWkBc1a2ij8KgN2FTjaIi3gT+6r0fJ68yKyE3ZVccbPbmQD5rE
aKp6E+DOjkqxAAjGEpiRb0N0qvzu/6hAd5Io7jdUiSV5HS0kM5Z05HXRtCuxdVuzxLy9+he0vK5E
uC5w8w2hLhiSZ/3H64J7ObZ1cC5b1J2xoPKFZ12EcSY+rKPpOSraHj+26QYVUD0Z1BMzXZrx3BKw
P08zHi1wUKkCIde2sF8cJeCVAdIQ+hYjDn2HvGXmRFZf69r/qgg80JUmPfuadPm4Vg+DVK2P3HTY
Tj+zt80C/fHfyF8mRrS18lnB2XhtZL84yoq8iu7iIeF9KdVykVAhPt1s1QJ+kvGT30d/p4O9nGR8
LwO2xls8152BcajRz4IStBqHDWJgRRSL3KWkBMSkWeQ52ezPpsaJz/XRo2jJJf0wyOHIdHc3rEPO
Ydrs6Z1PzPP4YegTCZgYYGAoVOGveO6BIyoi7z1lqW+yXVtOcpIIDRKxZ5UzcPeGXf38F1qCLxqj
EYwRIX/sKl+3Sy7KCSXTZL+Yizsl1ztN90zwUxQbqjjcRf3ybw5Pqx3yW5DM2I9PGHKKVJ+LUspz
M2ce0ruK6jcSgcR4q+/YB53xSD0U1QdYRIlDoSqUzSQJED1xb8cgcDVFCtSqeetyYkoesDYOol2Q
r+GBDRnYZlAfxaUgUINSqYjwBHAESewZUWI+9FVc2YieX3X+Heo2Xkoi23wgANSRbv0VD0YA4ehx
nQljXsXiPH73tnrWbrAAGzadOVYnkBJCp25DcIzB8Qr3nCHfoYZKuJuA5Q9owyyIfmdOfp5Vnmsi
cLKr30ho5RCflYh3bMZaEIOcWIAlYr0msXT0dH2bKw1K5c2stfH3Hi2eFld7yUSA69XxH9x8EjeR
/+/vFcMF81bDwHFL7I/V3yZQnU0MYCDaSU21vGMM72cV1/te9VVw+Ojjl55BtNs4Mv8Gc2f6yJ3M
zWf0H0++kMIuWBZi7CZftUq9Uz8GkLJKlyk5q63F7/T8gGoeH+URWw20gQq4q1knF6RtRjmwpyVD
rnCGJPbEHEkmDfEWWO+gThzeUYJQuX1Iv3PBTv/F1lvHcCnBcXzdOStxTMoLUGgqQeprHeCr7DbT
d1N/giDXXJMv62DIxFF/HVjaADLuzy11bncEC/Vk2TGNG2VYe9pzNpwMVPTuaA5JhKrzpuXViCh3
RFSZNtxUOO5HtM+JVSRIU9QmebDJjjq8J3J+3mGD78EvNn1lEM/5wjfPDT1Y0ezvHWbm13W/4WLL
s46tIB2zKLQF2abvgmJhNk9xyCJno3h6o6+4Lyc2K8L9TYVx+kglmJYUKyaNWBC2+y/ioE67/DQW
1DcTYwPIKOwmeZ1YN45BYAldPtFqjhFtv5s1P5O8+bbKn/A5Qd/73v2mP21HouKG10ypa2LrvkyJ
KFd+I3mPxYxZhFkKzPxs62aR1s2PqoWmXXvnGtSKKPHHm4Vc6i+5kLbKQ9gkmH+Kq1fxSGueEs4W
hSqr6MR5zd9fS07FzMmG4eDwFXnT5upgn33rbaXxu+r85OflaTIj8C59Z7srx9FTWd+jGg77ydW/
N0FoWNiKpXgMMJfMddZPWft+sDgrz1aKCvQ6qjZLMdNYcK6VcPfI68C76/iDd6H9L+TAvh9/m/hd
vfGcZ40O9gGGwpcWVYvd6V5CPbBLaBXz3PyCRnDg6vKRUKA4Wf8AIJIqx4GAaCF/Y2Fo81UX/QOR
ryjo6gsgP6nAjK5h8k8bGr/az4cuWavqmp4JONyf+5GfDD8ZmbrdcI9I+bIcAoix6iEhySARhSPt
f4salCOYq8wZ465yI4qx1dgFTPS/MBftGVzI5/LzfeEKJ8kRjv5ggDGRlvyQAWoV9B1DeaRDypie
oOJXRrNijLHLtsKG2GVbWyDVd8EG+/+qdUounFVZyy2Nxo3mJSDaKnnWuD/oi1u8ZjCEh7VN3iq2
yVg84u2HGjFDGwoquGFPXFIDveTbuUc5tWfvTfDPtzc0EApMP1ggpK8F0OVA52t0m2i3oBSXOA8T
Ld5XB1y2BaHKlSHobfNpF+DcDPSbzsOk0mXg7KoqoQzMWtoJSxrvSqWSY2dtjRSkYzS6VOPsEo5j
fP6UKlsTZcmLzBUJM2Ze2UmYsLhVmbZ1lLQBB76uo0a+ZWpwfqIjRXW4gnzch+F0GYE2IfqeixHk
ipWXaVp09tGKblHojsnktor1rQmG9QwdrAzpsCTK+ImW4JqGLsxwQRLYHRS6EZVkMQMGJ/5Ej/XE
fAVix94AQgdMTvRGC6isIzZ3XOJqk8l/0bB/X/xQ82gM7tP9xe2XHKs4cPHph7tCeHl6lOvkfHht
rYeA2xpi5VQIWtieVGd+6jzsfzC487rRlFZUjIDzTUahGwxFZDt+NHXnghGiU3Q/Bc1j07FpOcY3
gdgM6c+7mcWLoNG2lZmtSIvwc3KVNXd4cZXcXzYNShvYapKeN7FkWBbvQzPrwf1SrPC/kTUdW/FC
oyOk1VWzYEw3HiT+uPAkONWEQ6sNC88zGehPiCoSby8PdVyntAmb0SQvv5MCkGwosW/fb4TXI99V
LrbFljlzXWrzgcw6Ys9gBav48uUm+VNrWMBQ3QVs685eUfRWwikgA5f41IbjMez0iSb/du2htCbX
cCx5Q5peNCl2yUa3clL+4AxEcggU5C8oSPAxgoqz6jFOGSSIAYgZWITLaqUhlwq/zz6DABfWWjJG
lvqi4Vuy/dPPTnqv7zK5vM8/thKHaS4ZwFkTr1eFARb3se96HMxcBwUUS1OCENoyG5jlo+cGAOgB
+/mQuSSR9nURz/8ujahszKMYdd34QqSLtJXQdY969Psh4lnz5WDF55wsl8ScSrAfut1pUNWiHzlS
rqe0LFZdzejHuPLeKkSFhQrgpROGwUIy3y89QqFfCj8trSrY7jd3m2dQOjOv3+UGX9PtKrRCMAuu
glMjlp12INuLM2FSPGZDkLf3QA7BSsTOm+ADrjoaL7fKQ68fWEog7ZukcQycFZ26ShvYk9DrxdzV
oh4UhdXoe/XnlbbiDnXmiuT8ttsBUZ0ScmltizD+s6bRbo/y3Cmc6O9nZcUnforTITCodJECh5Kl
Jef3ucIL7RUW8UeRpYecnruKYEDBvhvWvFjhjc+PvTwmh5tpjmcpkMjaGuhVtzDlWxjAZjPJs6Qm
nBuatHBUo84quYdgR/clLQTAtB42udyJN+5RWq7JAyM8QteO4EUOoA6WlsG/9PBU3APoBwNnNEh4
S2GA4oyEKGk6oSn5+sqTatmQ5up1bJhrA6Ah19g0jr0Deyq34bry/GDOojVxByfaAOwYAQ6Rw08I
t0D3HReJ5YGlrKDarWjB1aLANajlSBM63n83wqP8ZRiE2aB04rgsUnZXu1e7vxyqB83FvhYGcR8X
C59MBbi+nMMN/UeheBSMPaiZVSu1TkTCsKMRDElhv1DT08BQLj7vfJhwouiIqJi59DSO7cYfAfJw
gBLJapLERYZu4e399AQ/J/Gy4sLORplYEqfg8TQVGqlEhR7GXkTHbzlPPuu+ebh7Qhl/7zV8bFQ2
Ntydrl3lBqkkJMmU5jR1Dz9+fajAGEADGKh05yHWtREiwZQIg3CE7rPqRX/V5qJJn9GFNYr4BOmw
eqoDnL9mYeqaTMMkd8BPou476F3jrnNvANAN3XxXnavABRzdJXGbECFMps81P9rJvGCbYCLtcXXH
Uu8w+u+bbq7P9V6pSFO/QI3s8lqtBPrGvitCviQFDcEdKFYR3tfo1ut+JKKy71SFYmQArPoV1njE
/nkf4OFvS6Czo7XbeccKBq1nWU/ZrFO1YyO7ZcJBNWd2ZRm6JJorTmayrA+U8JW+PpwxUE3PV7eq
OkIzbm96JRZoOU8HLHgRA0LjDkAbNt2Ov+NZEDEJL+S4KvKbCtT0xkWyOdh/Kz/su3hVUG6mV5jo
wtMmZBGb5/GyJIG66iuWyOysQIQ4DouSNZO+IEwETMOTcxFvGtdjHCCmbEw7i1Oe0ymSl2jqz/HS
+Xp/AZjknjiRwCDOA/6obfTTVvR2EyXbJEIK2q9fEbB71kV5lraJrV5MaX0zgWirStAtrhMoACuo
mDI6efeq+3s9IG/xA8XHqp9yB7hvCt5Ub4aO+Qsdz0NRBfMZoLKuuTsNJJPExhZh07D8b1uAYbX1
gdd800TXdtlNlGc8RFIm2644hGkiqHzobmKqCMBxVuTmKy8EXtnmGMwzUL2QoCLORZADP0C2IJ0A
ZpXl00ZlB+yFxcL1kb/tk/YXu8Nn+SGxKy43gbNphJZWdIXLXw02xrzDtXzlBfcYTD8tbhVfH8Al
JzmaHo4EUHx0znEM4CgJGfSR6nd8ca0Z039R91tQCQO8BoBV1EcZSKI+P5JPQUGVWizvBwwf13Ms
vTNq3WL8cATQyzeGU6R7PNttJQvaN5iknTj0vzblLeWAOeFKBM4OWf2vfzYOToQWM1sIHSeHdFTE
XiHpAPIm/ZL3iTroLdh8BcOdPfsEZxUkmh9S4zOrz4ut3ZUhaNuie7nSTGtq8E/XB3ZEY45kzirA
pLqYiAs1RozwuliwG8R8UIiu9srGu7/7yYBHZDSrhYm88j0iPqAgL7phaLGiCq/ULQA/HevYy/yT
rNlZtHOs2eXibdfB6uBaPIbPMtahMuLMm51qhRhjQy0EGtmyWyHcnnB++prvAlIfVMFoOIEvAxyJ
NUK/CjPFQiC9/2p1UWeXqi2K/zMVkbPP4M5lsugbFn1LbXd77ZNajA/27cgW3ANIQ43GWJse7vVY
7kgacfpg0h/hwMXeoZx+JB71krYjA9k5LjVtBM8H4rzd8ovbOa8YGQkyT8CwHicuisetnx0zW2EI
Afvv62j72JdWEV6e/CEf73gZb03pj5Qu8wmd6xCgkR4XzUZXo6A16iZQgQKWGJ2N49Z25RjOtauJ
Z0MSPpTZy2c0kEsDZkl0MoqOqJLUepm+Vi1em8PJOOQSl746dHCYaE0ZwhrlvQJheTlMaI6iC6Dk
PgK0ETNsLv8LFATqDIsiCyfIzKWh1KgMO6rtIHWpdtZoJKrx00dpdRgSj28qXYbv6Nj2E6x3pkAX
In6SXPcQymWM694cxsAXWt1zPYs+WMskbm17qNdGTdS7YhLfHF+0aQ0YLBSkbADtC/naQl8ggUJO
isD2YOKSLHfqc7QRnvY/1xNJcPMHXsZraRmjrpU6/YBhm9spqBIl6iOKt14suh6F5CHLOIItiozn
zBdl2Ms6B5zDyKpljZ2MpV3K0mQMeLfzRT3V7sYjrhoUWXSZppwddXlSaWclS/cuBnl+U+mdRUKF
EknhgqxZlXFEtXBiafv3Rj4JvlrTDNrwUtna6K7DROzfeyxrdnkDNBgwROcq+UKaXrM2rG0fCX06
uT3HJRM02ap7joYrowLCFbUvmQ5Z986ZtUDAfhfG6ODdQB05tMCEyWtDY2qcJFHY/Yv08e1AtaNO
EN5iw5wyie+urY+qaVXrwoZcoyU7AYwhSPLQcOaR8kyKhcNt8fvxCUQWi61YQjw397iVD/A7kco3
A9lMlbvx/2TZwe2q372WeiF4QnZtuonteB+bKTAyazWck5pZI104TxcwwB+nvkAIhAwJEntdNX2r
UjwB7rv5UZGOs0cPwocFE9gx6H7MlzocOlRh0TjdEVcGRtnzXyGo05sAnz/b+BHw68PGZ9g55Gnd
9wiihl3RCNdt5UhTmKixyI6lzc1rh29mycELyDneMK0ZA5R8wIdQZQnd8b23+9YulkEPnIBbX8o7
eIkbGPmK6Pp5DlfYmhNecdgUJlxmWrh5QChqai3ojcYrE7NvT0YfR19NrZP3ngebVWbUefv5ReiM
6EAD5ck3TDIxFk9XC+wFryP2PpKCWlHxXe65ug1ldx6S31Ki6CGkypOD9dp1IfJhqdmxpvK1ne4K
HCRV/WAfhQfjK0vG2y8Jt88aYm7x4YdHHuXHd4GqKgTENiUyzIxD2aU6BLf50whgrKu9WYN2d/bd
Az5MFJJXP9fEvXLMIkdujAlVROevVlbeG52KwPdTrZckTMi02Oj6o/ydMfEYg/EmQPAmM75VRcrF
SR0dle8n6/8FfcQnM8jCKIvMIhF9YbwphKuXN5+rPQ8wTCl++02eaOF4xE43CN6+IoSC9ky58qoy
uVfsNcyVmQJKCEb1p0qPpnv3o6pCysBpq3YTKS9qyQDcVmpnPh717eEh9UrqcRo/XmECZCvac5zl
iTrRjEmd0ofwC+gE8tdVQH01+RcZme9ItUhWG62IWdM7OKo6C/x3vqUbO7FvlW2gzxhC4THNEBew
P9OMA+jmUCtbFaS8bMeLcSMy2FsB+mngjrcqBq6mBSri6nBA6ZXscVgsMMeNS5Vt+iSRZdAfBj3B
KNdsT3sz/agORSOK+VcLZlSyWKq38eADG1KIuOdVxwHzQPC86quL5+fT49vcK6ARsTSdAKGtNZkU
f9WaWAgywi+XZmzHPkp040qdCMtyHorZ3v6CZUgh5yNl3ONl+oFPg1aBcNP7dOMJhURx8/fFGCmW
pvvIe3Hr15+4aE2h/LcGFzaNEXvakDh0S/BDTyinxQJ3nEsIhl+DY5VKyhm6FZUD2wMeKw13crJT
eF6LzG20mbM2w6W7gdFrVhPLbG/N89Uqku+Az92Oiik3JAetQnJfon+O+Kip6C2erXBjmYZz3uD1
KVuCh8MyIFy50JP74UTVI645ltyGt5Be3/V60LbRASwQCq9zlpNThjfYXbjNdOP4NHgVmLn1FPYl
WsHqfTF3RBZGTivEo3ykq0bCBjQFMSef6wJnfO43Ilq2+QRpQNNrs3m8RfFRNw1sN3MUAuWNwU7Z
2aS5hkgK4LdxJSBHa78HmBA/dna7m04lhBzXqHVUoBZm4y5XJn1fN8kwMYQUksfmDIefReZzuP3o
nYzhe2JlZz2Pj5VLLfE9Ne0qtO8/IzYbknpn+MBL/7s2LwDdVkt78Ai0gVPlXgDFeS4PBqvws5g4
B9pBDGfdEoo1i4Vj/cNEMhsJfytZW8FBoZwuegZ67Xlahia/eL30WUpWB8+jyLUu1ldyLZIZEfU5
WxxfFhxm5XGREu7XJUGGOW+y84pZojD8ANFezcSYG76SR3yzF6hOvnrnYSClHk06d0ti9aZxLF0L
T+OAQPz94SE+cHk07jpqSUuQDI/po4difRFIJtW6ImEkbATqQbVlaMDdNNB8GiNQrWmdUf6GLAJ7
Xxm2vkTxgTSxU+tvd2KQxy7M0HQRtAD3NKCTQIkCX182uVGIYmXn/qiZxT/OElZsQ40NcYQhBgt7
+bm0tRUQ4ALckeWNXF6j8Wt2yjgflw0cI89iZQtCKFyCN4Xd2K7dqpHfPpcSq4OZjXX1mV6igK0I
ixql8BFkBEzL6jaz7yj9SJIAd+Ir2eO9NCiQYAU9E7lsXLBJ9PnbaywiVYwsN0XixS/+GbLzV5z7
uluNU8c3PCM790Ez0MDYiYQ88woEYOhzCaz5HSTss7lGS8y1Mg0YJdE2PzQY64BK6k2m22h07Lrp
EIOfsISPnfVQoooBVGQD//6V8M3DL1oDc5LHNCko8IP9krQ7h7/qniixbmSq9ba7s/ftIWszVr//
+hZbBBvmwokmAA+NfIjFw7dni72tVPTCDT3qkXFhoXLtnCYx9V6VvLYL8YdtIOu8cPbq5QUxa5uq
M+Ykq1gKpZE0hc1Z2B5Fo/yk32b6Sp0C4YVs9B9fm/SFZOH3Me3advDEjaJkmmOUrWpBo7mi7Vez
v8G4xUnOIyl2XUHoUIgPuXRXIo3wjOQBeY5K+kNNT2yos6U5GJoq0vfE5fbcji2ZCbJaRbPDt9i2
XMdanG6B2klvSj+eqdBt++g0kwLdnvStdUIt1/qieF3G/Dp1YzMPvi1Rm6hzJjoFwrgLsXYgnHUa
FqPvjo5uA3+cd8nif9gHWsVpp838roBz5srQuhoB9RNpoHWLd5HH8EFfTgP58BdLihJI0assdbP6
isvRcDNBI/2GkpUZ87BL5KnDYZEsH4unw4xrrSwF5WGhToNxgAaj61jb4NEp4m6y4tyCVM0TwWjr
v0qSN5zbH2Ew285iggTclrFuxniSySDWYI6NNujQ1EkICGR9KeytjvITlbZjFnUE3lJtFm9r02JP
MtMhXKgpls9TPDsQ33cWRKw/ji/0ugd0khrwXsJcB1O8dZ8aFtbxiT1F3jZvC7BlWtpN1evf8OHJ
VAuaYzjFH0J3p2R1Zm9FkcUv5G7nxhqN+/vjiGFdZSqZV9v40NVtt8wURwVs7XGOBuvn3ygVq0Ol
lOEy9RQIaRNxA63VilLrsu78J4CEfz+nap8dlLM5OpcUhK+wSMP7iLJq5yl78do+FgHUo3SWTjgR
jcoLMFumEghmu7+SDHcdv5CNE0lgDq/hWgMeHp4oHqBDZ4X0ED5tzKbjDUhPL/coMayayocFwo7w
dfLRjROtD2bFj51Ww3fCeXeq/+ERG7ZMVFKWSgEptf3WB6el/PpjLGpCziT7OsvAyCA3zof7fXk0
WWCE2e445RquxfWACKPq/alriKZEfEIDq8voAuPgmpRdjo4vmnwQLXxZa8Im+oBBty5bqz9oBFat
xbX5H80NG8fBzg3YTSqXWOKbTDwXxC5X6u35G69gXJyvj8lOSqwq7jICvbw/9S5Vu019N3l91R7c
nMt0Dqd0mVxyNLypWtt/fgEH6f9d5KEhOPbOqkPvBF/1vBXT50Lf/qdPzGPo4YHe3kS1g7cci25I
HwgtMqE3eJiFYFpA+ysKCfwujPMssZKjN7AsPAP7ClXLmLX7vg3DuObgB3vO3sPSf0oOcHXFbShP
FkA76jndilhUBvp6O2PKEffcCT61JPH+m/XB1A+pQHScdaTpQuzubhZGwgu5voqKZrt2zb2b/OhI
f/t0mOboYlhE9NSp7G/+165NbuiDQT5/gGrKVExMrfUTSyJvn71r5i1zMQnFldHlbiNs/8pkGv5p
BySs+PdFjIIfdEPakxUX+JjbZNquAE1/NkXwUT68V6jHwdyXoGnggo0sq2nbp2CcMj2E3SSV9qnN
ilzOtFS09ossoRD8OTRs3mMiPDGF6mqfG4hk8DWRAjjJmB8nKmWf34gB33MX58Z4shdD+xixduis
ciZhyeloABFcKBxlg0T3MOxXfapnBv9SxNg93dWAnk2BrNfNp2cJQF+sKCy/YEh2ZULJiGOE4+Zl
M91BNpmSxNYJzvmCx4ra0D7yvKzymW3hNALT5zDl6x4JCpXsdqxuxqM59pQ5IXWTV4jJ3Okf4f1R
Wcl+GmzH52csOIhEWGyjFKEZLqRGd2PDahBF7tYY5/9cZ3B0l4/1Y5fgknQ7jtJppVgSp38MbkF6
GQoSR3u5zzNDdbzbrT/4F3S07VsivBYKAYuPBMZnMHVN5hSBtzfAOakBlUNaABYsQIu3OAC95ORq
F2+UdBl5oZXO6rc9k0y6Q58p0nCEokVFA7TK1dOcsE24xF/vcqb2Xf1Ow65nX/O4CMPA89UjHSzt
cSI/hhBmh7ph1deg6dzbLjurHJ8M0ovVuFOYDHCv/CDibZKjlWOd43+BJIb4QU5Z9JWEiE1qeEHm
i0V8A+tkIyVUP1WM2IBYd9TJL4KnHig/Qp6l2x2xWR0F8CUlcB2vQOHEFHQW44/pt3iEl3uivjw/
Wy1jYovb0cmmBxiBct4Yo4/CSKznRlUh2Gfyjs8yO9BCJNct3Ek25KgOf0GB5PDqSGqVoNXmnYAV
AEpDt9YXTI3lmelXImqg6qJUl65g5qY3d6Fxo7hgUZBpKhxcQBzre0XOaT/kJYy5J+8Ny9bEWMr+
xbFjW4c04agHkSJDoJ7i8QwJiHXEEejKmLP6rNgRuCrlaGGFzmbUHscNdoxVidryWX/MIMJ0WkEP
FkpOMn8TMHQ/jB87575khF0eBtF9a36p+KKo1SUyA0LMtHXjdF1OqkA/xVpRH3RcHzrzXlcv8cvF
NTFgYOXRMZYxMY5iSaWjka/6/mD2YMdCkU3FBStFt9AMbP6U+TG9fjpAYjGVm14e2zmuPJZhZuAp
XaiQKGbVS/ld9UHHsGS2Jyy5MzM/dV1C03BEH7xql97Nztww+fxiQ4jQ0Zfh6EMfdi133iYFK38D
9catAUWs6uW9FfR95cbZjwNb05+xE41NqYSNlyj77q70tnIM3/P2JrDlDQrxq9Z03BR+sMAJ2eT8
6NMnlYw/+Mk4njHUK+TAhitYsdIik0yKjo4Sv43kx8OGn350dmSlpCoCU/BiJee5P8K/J/O5Espo
JEjCoCpxbgo/2J1S3jGisDahxPHwxl52YJcnLBEeLCzD7YMUi8e0NrXW2LSPz9gWrnclszIEq/ij
LW7DiHzjoM8495TTI1cUkZ3heTtipD8tupIepDufqXuwZvVCyA4Sm0hu7JCmuBD2/Fcs5kUZlo9p
9QiMqFcfIkMaHN3madq4a657vZTCYSESDEJOzgol/pqqLfpRCGF3BiPv6DFilhcJ4pmhowuMc4Hv
VJgKwkzHp9c+ov40XvbDOY6T48tYMaLKjxXr1kkCNgcCKSAfcrS2cZ4uImCfOLmnCWV3PS3Cx6VN
5YyWOpgTOfb4p1r3MpLpQg+20A2cGeNJoqZdc/dRsRYbpcPWbbZ6uuugdAIqHwVWdTIvKg23hW8C
ycd1yh1MboorJESkmmGsNLVa4gC0KBGSyOrpNNOupUFSSAwG4zPQZ+q9B8Y0pHMgMtK9jUT9yANJ
6YprNbT1bAAQn4pI0SaF92pAsdfeYnoCcvHToACqkj/pklnwKfEVYzplbzjmCKBEvzkRxqnoS7Fl
YpVg7obCG2vJ8Xflfuwi9lpbngrcp3r0uDQxOVOQjunQW/kJHqbSXKsFd4nymY2+0v4s1py7kJdY
Zhi5CbJSjrhfEeLwSI/K6mUQ/zTkabJQUfgoJpGMPr6O6joW5gQjtN+4ZPU7NfjaOITVw3I7fUDa
E5L8g/A7jcnn4LL36Nv+hQs24EOhcOuSxINWHc46o0LkUUEFw9ms6kyBDJwr7oncbfBu1rn021Sk
xkw2T09RV7I8vzoDG+hfAVYSA/8mkPLtu0ZMYznzh4e5wIpCbsrEJtJ4jE6OM+VAcpW3qpqw0TOX
SS0dYdP5khw2xohQmZHavQcQnky0YbglAK/WqPAYl/nb6GdnsHiCO2RoZzRvjwvESmu3ClfvagJf
AlmE6UcBHlwlT06Cya5XDuKPcZfzUICVi85LsXbFhBh36UsmVvq83Fy1k4I5iXy3gj589yAJay3r
DpIJmRULY/SXVzT7vvRMfVPCV2ablp581lbezLlXXX4GF4tVMcji5Y+OVAjL20IdJjD6+BdvGsUs
IDIVFKU4isZ4BwSJHt7LHOkGAzZfbFU0thXB7KY4gwLiDKFvq+R+L5oFR1H/0Zw8G67BdlzyQGS/
fDVBeAX6DICVOMiTs+6SxKqo9HkSfruplebOgzGmgF80oqkt3UtyEcQoeaQC8I7yG5BDFZcmF+sW
9fttsugyuVnFy5Apx0rkGxsnMtXHWOhG5itghWw7HAj4j+SHw64rXfgneONR1AAm389oeZWN+gWa
nmK0m+EsLlptjXblujtp2GU68+4VOrFnDISYxQYrnlk51VmQLL9HbwgEVkqfeo2YsUDG9MFUqQBv
2bcnUwAUYYlrkAaAi4LOea45euMeG1v1LbQzdKWL7MYItinDBOG5wyHZgna96Y3JgWEtPZbi0NO8
2Mvv2WQu9LUEb/viWxxMQjtEtkSiViXlhAoEoq1lvrtNLgdOLOVvPZ7TaEtKg+0rsBmSpOhxldk3
mdj+qShfy0ssKqsS3J+1YPxshK54XUFtMUoJuLWiY1qYPpObr51eD1SvhMm40WuyLVb2w5646pGF
YqGZmIEfa3jn5FMgwfkj5XtPckmySKMeM1vJAtRybTlbNNeOwZIUl64ICAVqoXfwbYGilKKOo62O
yKPriCnTtSuPrbfd6rd+sQb9Oke2S4/R8L1DFPR7PSbktrmDtQqR0sOo/LUI45kKGS8LrNg0ToSu
w8gs6wjtHgvYTGXPyBvTCBpqUlNUWG78FP8sHyMt6gSg/5nJla3rKBTB22dIHMKlJHN0PKrcuMHN
nnJRDSscdfkBnEDiaajkiNgQ5zatLSN6QNc5aF3QEOAZ3DVIoO7uH4JgplgadikMB0xHUZBp5FrN
Hr4OeeM5JQz7zQnE4ZR5Okswyi3QaR08cSRbC4NetE82HlHj+bztF1IKko+Izc1KmqMEzluYJzdO
PGxBeFvoQ3gfpYXnlE/Me0FIJvvTDqoggp7gOxvat1h06sQZfO6hway3luC7T+EOYPbXb0mejx40
jlh7ysodVKmWVh2s9AaJ1w+ax/Fg54Ed/FQia6HGlW5RL15VJFI7MsXUB8gVIGsaiWiDBsugvBbN
TqcR5NngCDXjyF0ZIUq9ZZTpQ+OhBcOwiVNbim3yXC4yzW7vUkeL+JqPZqh3iCkJpk1aFW6/uCmZ
lZJvBspNUwL4/VYlLFDG6osgo7p7WydDgJFQUSoqBaAXTB3W53bgoVMTQoGDlojCd8A2k0uzMSin
0+QVuTpw/DtNDBdy69msR/KAHZJTlbCPp9VLCk0LRQcJ6Tiq7QRNoPj9HCUv3H6HwEzkmH0UWXAx
FWpfcpehzHa4Amf4oWEy1vAW9Q/6/XOOrvH71CgGLITRUSmO2joLhiJC8MxBQO4bW44NxzUstYSw
NNPf129K6ZIW3enRzoiz7XAWOpH2drzd8yy4GOWv3ig1xzRhueMtrsyXuOR8n/BMepL+myaUpNwI
Mq8dM/dI5XTnKkC9/F2/p9/rv6INEZuesIXpzqSWJHPBhV1lhmOwbGxCGBnFyVXjsSArobJe/U1x
A++twUMt4/j4ymTxpN2mTF7uTsOvIkL8hpydWLxJX7++RFmqSGcg5KS4tc0keO5yK/PQ4tRDidyJ
HdWE6ggCFdd/UHkLgmH0bHF3YStLIRsiaWjFbHKx3Jmg6A57cN3CEG3Q+MYwAK1F8M5udRY9BgdI
ADN72/5uUeCFCtxp6mHEPe7ix+EVXqEvIwm4kWKjIgWBfT2vCNk/fRrY7EQKf98AJUP7n8Z7OR2A
TO1UsT9IUJBDrbSnUfpWt8LNm+58Xou71BolP86f4lATvhpCtAaQLKtJ7vO4EuW4TdMcOiBKe2s7
aO3TgnmgCSm2N2xwoDzAu9FxJxhIzHcS33/QcXhSfEZkbIe8tvkvYfZMTwcS0mVytlAJ+LfGrUg1
aBuBkqwwJXoS/e4C4eP5ZhBBVT4+C+jbC3nuRZ5u1dAEdyFqgSWBAeawPInq6g5ZrspafvWQJ7G+
fla2MlGGwIhXAAiCXB1+OGXnEd03C6V/kO+PTJRRLENrH7JJVmMMFzRPZPho/8G6inPWgwKujTlG
BVrSM6Sydb6kQHfGENyGQ3wvg476HzzBr6RQ9ANRebX3rfDtQHmYOfj7Gsxa9oux5bexGsIlN15W
kIiQtXhoIfYSFchZkNrO7TfArMXew3Hji8fdhL/HwtBsuQSMpH27s3MrjVWHBsxRANqnrMAMnLAg
c/9FSG1CiamOeBUcHyQERS8IEW6xjDeRFVSTVEXfJ0ggdBnOAVaAFO3GT5hVye3e2w8BlZKRhbS9
3FyFmVmz2hOGk7o5HI/cWPOKNVMPUsHWZe/uqLix29Pr1GlGpt1KFJDS1sFhkma1jMrK0W2HsXhS
Wu1ON9VencK0HRHPFdZjcUqpcTefFPeE1bG+m0IT5wNqfy8A0suiufJE4WWBLSwHT75/suqShvLE
tCzrMcfOqOBo88zicgbXucTxMtH53E4kj/O9RN93J8ls8/J8Vsvy8DpHnUSCJKfMRUb0vKdsaM0o
rHiJ+XLLUz/83o9TfzyAP8KPbtjxjfL1Q0VPInhck9XTdXqH18vv6LAMDDyTc8fyr8485DmkXFqi
fzt2y+LhXraWSh6rXSwQ95kIKl3hvy28QgCqAmuHzE9GnlABDVTJ4NE6YNxhVEa2B2UTxbu0/Q/v
Auej05/n+/vzuas1H3E0Dn53yaWMtua9wOJfIqzLu2LBTVDEzjTMEC62AuXhinN0lEqQAMmxYIFO
acZFIBL9jKs9W46Rzw+Qre8goWowEkm9/3wVBpv+Itan9n/igAK50s24K1Y2QXb6dgxx8RkjK2ub
zWXeqvjmWZ5insBqK6SCxlCHBkVms8iYYKvOtq2/LnpeHfd85ZoNG4BP8+cbTv7itBBaSb2g+NVP
efn20P4dI0QpQBvH5s1MCtqEuhgNqxH+OQAA7PyiCNwfagz6voWTOLId2TX0Ix0lR6j4UPgL905f
Vpmi5EBbrbgS0rsGshlXfzdFxn1u3PLmaDM1lt3w0M8Vbq1y2yXUsuE1AD9dI+cNYgRZ6LK8VMxL
nBQIhQnItnOwbPhF0zhaeOaVZF4Tk1zC9m/lK7aXW0lf7v49rywUAgEipSit/TgnvGbwc9X4v2y4
2c9OtBrIYfqMGMNYO4d7oHfdOmS2gO34qG+dklpjk0BdNiUlLp7gEa39KzyhA1OY82ePtIlQpXpA
RHkjx3OhimAypaFtEhUVx5zagSMcLz8k7VNEc20kGZp5pO6MyjuULSOf2nx4vNZXOQ5XefI3fZHL
BYy4ewYXqrYQK1NQkzgwvgtnKe1tDf6PeREZaErUc6i/W8lVM4YQJbwPkzMAjq0APqLjZddIySN/
QsW6DH6oqOacvcn3rTX2KgKvia9VYGoKfCHwxyaQFYhipEQnHSRL6EdwMbHTqEEJS7/YPaQgFI0u
hsHAyAeKoGJvsqJgySbroe2k0YyRftViAOOsSyDko+URK7KKA2uDv1ynriKyaN/2tUemiwgoIv7l
mne5YGUu5cfWqBCoqPY94THZi/21+ENkE0660jdDwdseUTn16O7gFbvGFnpI/iMfiu5pbGxArBIY
R2tdziuridp1WtT5hP7whEfa5/D933iJvM2Y0gbAJlv8pba0KxQflK38WilA5XvoxLh6QLe8ebq4
J/cuDCL+2yGJlxWmwHxzSAaiOf28eyz2TVpu9g6kUHs8+XAZx+fANaXreojBhzsiBTDT2XH2lCEs
byol9jBZ9CsNRU5dZhXpnlmaDj32yWFo1wTXlgIy4brv1Miwf8I8lYoEbyd6xIZ4SxFF435cWY4R
6p4yd8sYKBw4TIQgxS6l0A+b/6DN8WUhsnnPScE9dTdXh8yeTzHBXJtjZE+bgTcB6/UAs2XKV6Va
RUN5b7cY9my97pes4e287deWdURg8iN8536wq6qnillTMHZcF/6pkD2cMUEObE7r984lrZxheQdD
KxK3wLy3ngQRJW+m1P/g0LMzmod+tBtEVx6vk1UezFnbmr9kUD66N1Ce6J5D8SBsNm0KPuNmyNlp
sbq+Rd8grdGB8NqRDi0vwM8jLUa5Cx+SnlGHDUi40LHnKN3MoPnKzlrPcClpOz2GsGo7Q376sAAY
/bltPZJvdlr9SKP7c//fHtSb9eCCQEc6ZNYY0KrSYXojLOrYA019hdVDehS0jGrvElYMm2tZfeK3
Xyi+ht/GlBKluyb6mcG9UTrkBehBrSN80gblLZICcoEFIcSILvpTJKA4AFw8Cd6LTNAmgp4fXCST
ulgDvqqidI0MjlrKdqcZHtScnuCgQWQYJkon2UgF1O1DWMgPIOHI+kgscp9Frpq9Dxn/Ov/YfWJB
Nzyp8v4IJjDVV13oYZG5WmxAzg82A+T99PW5EYUShx2e57D4/Kg+8nG5TqxcOPNkoQFpNpw7RPv8
LbciqyC0GpHdxBJPAVPSqVGsR/++hfIINfHtlrDKEk/4cpWkEQq/oz45PPsr8kuA/UirmHLtsPO0
lxwaJwYgYaafqVkT953hXqfnmcQ+pXSi/bEuV7Mc3ylbPbeHclCbK1NwTwPgMfMcP5tx/yGoOeH3
9yNhpJ1VXzTJDvL0Ev9334vEjvUUokupmyoipth3iUF4xvrHGnvszRZoI3AggMAK0uc1TWlUgauP
4pS7Bh/jMEvYxdcJxBJNQ6UXbwVdbQjGvMbauL7xsig1gNegqnvZg2iPzikPW5MyYk8d+GeNpuCz
FMzqlojshiGDaSMqLPIi6zWWRFKnFpJW9eava0JcbE25fwEVRY8EIXZDJ4x36AU9fatDcuwu+fAI
IWrxGT5wu7qD51eehbdmdof+bY4Kbwsf9hhhN2nERzz/jEivG5E7/NaSsGvoE40lz0A/J7eDx/02
DB67f9vZ6pJ2QMLEsgb9NnBYXrPK+2eU4V7FPEOtlCeglWda0WWjodugSDc76vNFrjuPLUEV4vMF
sGqTc3+x+LPJz4aqWFyC6uOSHc4lC26ycuQiY88aaMBzeQK8LHniT2+kfwuMP3oko64HkdvvtzuJ
f2MvSZW235ZwP0lmhSsJqCxn1Hhubx0z6uOQ9zeHuZC/89XhW83SbgXvAf4Cgo8q4eZDYJ6RsTt3
RHVU/8Fpcb93Wi7IZ5MuMqWU2p6AuAUBr6KXXRQRTSiPEys3miKn+QNILskO7TOztittZvUrLjUA
EJtorM5h7o0l61s3K+sO9zaDWS+pKPIY8U4KwTjXY8jGVqm4eUW+HdC4NPwYnEadm/2s5ucXPI/2
DMVUSlS0VvZxgT7F29ofKuahWCvN3LXCWvmxp3yjSL8TXlK+716usPqCDWyLZ2NCOY7jFjR6XlJl
tNzs34p6jPXuOdf9EVGAh6/lY3zcLjKECbDT20/L+hJEhOPykrbPLQ+FKoVTB9glLvzGtqUC0Z5T
2dj1xNK15/70kOwpGzWHVWctpUFieZqIdezPtf+jpdN4jwkPEQAyNiqjdoKtGYvhlKP1LoQl4PQX
iVk2PmfylkOZtUeeOfoewN0Ad8Trel52m9VNgF6O18QbrjLKzeXhRVe85XdBsE44BXBncXTwWRZR
8Jx6vQnH9GkG0CHoxp/YsU7WvdsegaO+u3drITjrWqR288v0PEktbO8nKEjgLZOVZE9V43YbX/dG
wg5+sipvpl5WiiY00gSWqH9IPyYO9wicjZFz+p1zBTyW4ecMUHADgrCNlNa3bJ12qcnutw597Ds0
9lSYhVtNNKbjYMa+WpRMctOEwrnoHD1xO678qrdnMC+w2tyOAQB2wtiYtx+Sni/PwfobSSc79YQl
KLNyxd9kDuOywIzIZ6YGNpljnx4TtiztjlRwcUbYvsyukx9lG/i+DwBt1Y2e79VilUXRw3JTUUOR
izf1kmlFKwxmbeglxsBPH/5pDmKXp6FVp70lXKs5hknhfQ7iSc+aoJJwuWb7SlMK6IzD7oMjjDgT
VZKn8JnylfwLF4hHLKHdnYJwVDSB8CTUJTDS3RG0Ta1WcLTkmDAdeNu32eDjqdZbL0koqjr/LTRB
ryJk02Mfkn+7hDW1gghS4ChmcBkVEbi8+E3T5uhmgEMhxVfWcHavjEvSCdYuxVEtgpz3Wg8LrrbJ
0QanyZbKeY/ecc/J62+FMtP/rTUCWGHNqz7fgt2gnDt2cqSnRYeWdHdE0/mN9p+utBagzfWPCE+T
1iSe3ztX+zhC42UHPrBEPT+wGIJ29pgDglmy7hwF0LRcm9JgCv1Js4qrS5jafDdUwQr/mQLoBVRm
Pzr2y55/PHSxE+SeRtPwtC+7NYKCiOfq03HGvomyT5rlzbDD7Y2Yl8pCTesqmrYI2u8tJXPwSSMx
zVaxRyY6mFiRhFr9rfC+02G3sREELCzeJasV/149DCbizJoGrzV2d0ww38q4SrcYmpQb/5CygpV4
koZFrWy4cDJ+K6jIofQwmRFtGbjAMXJwvmQjIK4UB4fBvxqnjcl9Pv27RUb5izpFNbsGQ7T9vxvH
eZnUSM57a4IcziyaGCcAnBCMFl8qNulipf2eGviByHQ6qKHbmiCYDaYSzoJsaU4sWhyoje6IMF2i
0Yys15ixYGnvMLz7nwfIu3XaKnI9QFdrjhiKofX53eahARCewG+IgXqZsPnbO+Ll4dffYIT5Bz6y
lzWxOI8v2OeGS5jvuGiylkhbphOJs9GNCKKz0kzTKBxP8ecOJrqiganaEITK4mC3zZqIgmgEJjvi
ONuW6GsEta+F+yKp50l9rL3anTDDEs7PsTUZP6u1yh+YtosuzVPvru23aGrHe2c0f+/rlfoF1+aQ
nA3lRPFdwstH9MTMilWEhk6QRLLW9tkMtlOPfsY0StyRsaRQiXqwH/STBSKHAgxVeTBvvkpePjL/
eXlz65n+Qu5RNfPbCuVhQwwKIy5PtvJyU4YTDQrh15LcMOAqOJ9cFvjYPXv8eAl28tIawKFYP0cC
V7CaT7uwHNNF3AD5itfaMMwdHu2IxK3JxU4Jh/C2yQcckkMmQqzYhaIrY5gKNtLEXXxM+9wsnPqK
uBZDJ+a4BiZAQ+M3bc8/NTbO1w2+Q2HuVkrUGKrDCiXp/s/N7VcOukklb+EvjQDFh9lHugr+CGbf
YOC9UU4a60WMiAAyD98PlmUMORvI2kkIyzVjOTmnICIh3ua19kYDQqott5pGFvoeNiIan89x9I8l
2WIpKfFJ5p2XnnpWVVr1otD9jnIZWDzL5LtupR1XFibaLKuSFFjYSlPg9YdZ8XgVnGvuUOijnMTy
vVTTLAj4jOOzFfTmHYCxu9EJywUgCUFZmE87wqaFV/mulWI/xUKq5Ue1WOYGP7C8+5P2WuOhcJUj
2onC2aX4wf1HNWapEuPw+CoNdRBpsfhd83qq/haC8ZQtBz1ZzVHWgCqRpJf28sEDMIgKvvcYxeF4
Jz1O2nBFKNsGMBtAkxu1QjtYxvH/LHdpKFdFWEpQBZXGVpFuwJzCQUHk7EmzJElx+FF9kEI0zVdJ
PibT65dEzaEgpjrHjHc68yLOV5hf8yaClUVVWHO9vlIo+gVDhP60l7UFt8Q/hgPLmvpItQ9ceX+n
Yk/NKh+eriM/fQAmcMlYmOdMSI/HLS5XfWfIX/xzaIWMHlCT1IQXVdY8HIW04s+3T7xvjEwLKLx0
91RB4TehHJdUJNdejVyPmHKrG2az7l8rQeMIeCEw+qoK4Zj5m7txj7okcDhoq/layYET43YL58cD
ONajYpMxgDY79XXJQcAXIzhUcFISxJwG4hiNEd2G5Z63GkVkoNom6FcK0YIHNotUxttWfoVt2TO+
YbL0d1SbXeDkRKTt0cm29e4wClu+qGU6IhoUDEN7BWoP3wEBX26wTxjTL7aGEV9yZjuA7b3g3xJX
sDmjbvVW0m5cxo8vAR0quxAYQVnkNNLw3k8dwNr2F/jHvMTcsWkPXeGlv2NFPik3Egx+D2xsM5DY
Cc7FHKv12AU9g+gBIk6Jl3MZh/kH9jVr/iOP+TEAh+qC2r8IWnzxVC8a7boz3Vlkbpn1XmNAbGFB
Ie3eVvcn+NMw0yxyaX5gsH8L8O28tN2TP68V941ElM/nljBtKk/KNspOSA2Mh3HC6tMc95iWQTh9
1CJlQr3KSeng+DsE+zITTIoC2GO/TLhW++say7RP9HDP2za6+aedn0dKDC6O7xdER8iVpfu36sJP
DPt7dIHECozDL59NMiGzWlppgEOhtOw0KPRXf+Mv/xIynD/B9S51BAyWifdJz62qaP6HubeGiNG9
LnWgXGQHf/ZAZeEOvrAVU4l7WNTWXPp9xmCekatuDpf7r7zzTOLf1JSOUE9U3vG7SRBzGFbPCbER
URqA4jXFYTJhWulL+6AEPl7zdfpPrt/Z7GZm9GcnswlN96lFZ5UFeV9kHrqfN4S9aEyrhgC2MJZ3
7mCVWuShBJUh7nFk2HMRKpI3YzN4jQ69osnfdDK1g45FVgTTyTT+8RcsjgF9/m8wDjBP/rLQjOno
AxpBygdvRbbb59G/b25UeHbTHDKth2O9z+tS7F1UvbuaO3Eaj6TxhI+I97AZoNYkT7H8BcjVHkVW
+J5rO6urpBTZ7n+eQe+G3pxc3zPeBkG2ZwUHUD128ZIk0OtGuq7QR9xGBxWgcaFDefkmkzHb8BtC
dMzaVu+3O8XwYQn1SMef6o9mNsaALAFWmRdqBGetSOLjyn3v/3bpt0NItGjYIsDCYFFLEHaLp1lG
YQ0CUG1HeKSQLEl6SUmtmLanERgwE2OnLtxxRBVZbxxokVTHkVIE8R+E1I26Un6LybWS82r4kV1W
/+71HMILs1/gjavmWvkxkfwefTBTnO4SAdSLV8TMxReo+8N6nml6nDcJ+5UELER58GUfU+VMiJOF
+KKFhJc3yhFT8LycAp7XVhDSwRfnGzrv1fj9zsNxKvUGqPZMCN8XTfaBrTXGpJBJ16uy2IxFX8MR
4tC27QBfbPhdBXAhrV1yAnJorcR+EJagpZ+NMWWgMn+JZSD3/A13VDjig5xWM9J5xlPRxYGZrBqD
R7zmzLdjM2D5PUpUTNXBTjRMARtGvXMPhJSJ3e4QGEyKAtPlhw5Svu0oAfcXvAKivp+teHcNEp9x
taaJyidoI27M0z0gFKif4yc4EfL8TOg5Y3bAlbiX6obAFMJ3z7KEM7aygPFkViEZ4CzR16a6TXUX
cqBbf2DgRfu58JDr9NVODkC4iYNH+sv/EWRH8+2GG84LRqjx2VkH0XFGgwa7hRvXf6K52Q40Gxka
4OgDR/lbKRReFe4dof8vDfMxQGUFZam0egiMVkrxxJsZ9NgxwgH2RRgDMdOvHb6zQCPctMpFqeOX
EXVVM7eYnR6tEVyQViafCVnVFy/PEzuq49RGWrV3cgpERChHAV/CjEOjuM2H4VhKqZ1dM21mW6vp
AOHPtk3vSWtrm/2FuOy82mBFoi/uSTLp2GKL2YkGuDt5tFgrhsP+JWkKDCyufcdC5aTjy0T4TA2W
6kspGK0GWIXcbhA8osBJKbE5j7WDna7SOwKjpoU/iXVz2+L+4pVWzFgvI/RoiYbWqbPv+k3GZSiI
9U9QbymwxG4cnjomk8FBD1wvxxxcQxISgL1mitFg0vfipah4jzRxW5LP8p/LVntPG1+zaXhVUDgz
06VqKFshY9sdLyMT6yLPnHkj/2ni5f6JV9xDAhSPNPLFsb3mQZprJ3mpxVjlNUMHJ1x2ZQHXRB++
/wda/vSGrTLtXMm1/2ctrEHYUKXoFSje5DqaVA7R4nEC3z4/pde9MKkUxP6ecBsADdN7Buvho3Ma
i+AahAYgiI8LZA5lrqXngLbaGzOqgDR3RLBwm1cAvu+NcSzZ128G95O5YpYBQpz6bAqkjj5piUvt
uYEmSP10UgHeoDcxzvSwKfhWjQUhxv+ql3486pwZXBqUQY5dcpxTxMVZAHToNh35iAES3P8VXc3l
xivQYJrp2UiXBGA6fVuGJSc/IcwL+KWOlryLj0MFM1cAdQdhFZeVKyo2OT5YK3Fnb35sTnG1CMWe
FQMth0ljfUhA3Z7vQx3jxOlF4fEMLpGJg9kc8OQspHVyIb7asW2HaHt9N3GGtqzJjAuYEIAmdbvy
a2a7OmOVF0acVRGQFEIcyCbVEGEzMe4213vadTdw44JZB+P6FgSOkEXM3lDBQQepE8fzSEMiEnj3
TX6tcisoVoStDCREZvu4U8e5I2vqppiDwAIv275eEs97yslDX3Ln6VISwP8EwA08oyspP+4hSNS3
A67o2OdM2vJUnnS5GRugm3+Wh49HQ+dmKDnoWGDFHbA/d1+fFcj6Nt/PLnosEgXINRl5OpLsOwLj
I0k0CrBF3nnteKrbQe2heaqzOqMgDNQEW7HzzHxtCDdQB3ToE+jQpfZKh09tBqo2VAqNgPrNspSx
uT5j2hUP8JN6Opw3kDHfSo7HInEmIhQ+DGYNG6xD3sKyrjuTh2vG90KY/ony9dfEV30PjPKgrIZ0
YLWHZbD0tQvBDkot4con9MMTzLZEzDyq718OLIXVBP5nqxMGHk/egJ/7rFYZM2JA2HRsVo+KPFnf
IBAUrWUHz4k3prhPbGqqApq000IQ0Sh1wO2ddY3FF0EEGzNNzNC5N8NfsSl8rcxkR9d/1/kJP60s
Ox25TSGgrsm48K/ZrjYNJ1sgQ0Zfznqmn7m1WYiA5vrbgvnykLM76Q2NQCvgJZ3a5HurxFFjNlp/
vP5B8ptfWwIqBOPBnuWu5csLp2lC+NrLscoL01e4RYdY5JkiFHxNOnK0OZidbXW1svl+njJPrnoc
UhIcvQL8YYoS4AeJ31drwsMJXSGb4rSsvcVrIcnVReOSkDi2huc8VBqj/2yPiaIwootZb82AtAgY
KX4xpJwEDefY2tVo2as8ZNehr/3ZY6bSA6nMDIaRjOamM0LUQ/HjnoVD+vN7w4BsI5BluUzTuAsu
m88Pm1m2SRmbsca4X9hjYgxlt1E1Mr9HH0z22JQPDTcTr7ERbj/6YaqmMWT+LvWLyVGN95k/opfg
QBMaFoFQMy9UUbFl3uOaMcUSwOGYBBueQMULyL5B/xWT1Hrsa92/6ir8HkFF+5Mmy8OStYkx/2Uo
P5lA4diNCfBPCm+nYZxYdlhxLOMcP2P3MHN8TBc1zEzg0aKYYPCNJZdBq3l+LnuuCTPXu/Y/xZ0j
dDd4uGgrD5CbUBnplo7AdAFw10w7gE50a4JyVjXJ4taKEnFfv74v6pAAinhYrYpqJCMSn/SpmuJa
fscgC/YciuURif/oRppWZ5NxDAUQbxomJTsyJ8Yz+xqIA4RN/9PSNoVVpVKTdQOcunlPexIU47G1
3ZWac8gNusj7+GZPXuAiKwsQiM2ntz1hbLDxvYjfT3nZ0NmHEdlWKJZxYpUANsLxxjeI+dSrHfvj
XlDS0UfddJZ7gbOK0A/aEvYKIdUqJ3GQnJWoqH+jqixx2ptE6yri5qm2RNPIgJ3JU7w0tC6TpQOm
nzDY5EmBiY/O7O8lSJXTU2PR3Oa9ehUHfTZUV5UMntSv347K7WJVEkCMSpr7Ry2l12BmEERtcgy4
O5SxYcu+4igU9yYZ4/gS3gdE0DBtncGCKVLvK2lKZv9vvTwJhF51t0mUm89Y+0Y+F+ySBAFiADP3
Wkfn4N+VBVCKQGUCvnoyTzt++oJEart3DiEIAYgzJ1FBr9U4lxn53/8KqgE8IdfRLnJPtTfS878Q
IvRcE90IEPnp78FQrImNh0GCjOtAsz2wMjHDP+ZDKCN43Qw40S51myksImokwjfI6QZiPBDCvzPv
MPsgKaXtZKZVVbilLxpT/xHCud6/4Vsvvt1vA4V3+WfqS479+QIzrqeriN1YZ2EkY5QdiUNPI4db
2Yyc0OD0xDtTULkB4S+JK3Di0oC+Ye8ocXpwxbecvByt7bILBy5XKX1Z78iGnU8OgAtdrrTVACFb
a+QjKqCuZfr7pGBcA7JkbD6SuA06ifITsXNR7EkxpKxJ99/cp+kOZbjoEgIctBax2QsWhZUO8iQk
qnH57LnaBvIB+egG7zvtMsWtNc+mMSTrSc2d0UPYjS78dmxdx0PtWpiyRIs6ntvSFplN4UymdqNg
LI9OUKBi/HJJY3NZdC9HX6yiT7yDK5Sl02At3vdzOfvao5RVgUfVcbKyskze9ZcPD2XkCmmdRgH5
FIrzdQkcYiWLkuUYKZ0tgbZVFwKPtX9/wYfMs/6Tqi3qKitMlz41PJ+cfpKUPI0+JpWJIYgj3gyN
/rb2tm8TAvHAGmL8Ehi2DoAOSpfFBjkbUZYz2MueJPy8Gw1H8yTbxVBrAXvF/KfzUJj2MYtu3q8L
ar+OHFj4yyuSjgsE6YyO6Db0M8f1lsfgYCq3GzfoN/O4ybeYA9rmalUu7cGlLGlEw0DZ9Z1jYvkO
PFhNVgwcxwzRWE14iO5Opea0oV2bzO0BsWExEQKvnf+jGrY75eBsAXxDTuI/DtZl0xphWph9iezB
gf63AXZhx2PIJN1MoFZ10O6lwf3rrF3yJryt3quhYrqxBny1VbyxmyajOkZtFHfE407Ajc9HcGKX
TUqquFfu6zhgck/Z3uSHk0QnJf0WMhfiKC3GjGQGsQ0T4z4+/HCZRo1SlJ+ApbDfz6BYI10bwCxl
TARa8OOAap/8e2yv7pTQFVO2plzbP6OYg8sU4ksJYxGrXyK9Gn7nsW1QfIRMAh3V5CxhT90tkFj1
Fxe4coN8f7AeSYH+vyFMSAPRS3S/7tPzMbleOgHyl/Iwcmplm0WqjMMAhCOrCltqNyWcb/8AzU6B
HLlna4Sp8PGd4wg6xAzlNzoEvJJLByHlgmXQUfWvbJmAsouQwDIy6ta2keXRB4rZXA8Mhdm5Qj6Z
HF2RfMzxGxp6I91s0wdaswnZ1x3fKU0VgTLt1aUYegC0m/V8D4TdhK+xrxmetMtzizFHhNhF1IME
7sQKjYAgLJAXWExHKMKaNZuSRRqOF0lG3nSfxdtsXrF1/Xn10HSbgqj4q912EwYHu2uam5QxwMc+
qaHK+jMW/eL4e3Cj47lvPOXosegGvTtajHMzUX/+RypYL/bilUgjnTvp3lgKDEWkzwS/UiOGVihW
gcrB2g5JBpy/GSeNLONlSVFhzxNz6pLESjcx1j0tpVrhRNdyqPPOXw5E9dcGmDUXo99f9GqSGox7
n8RbP2AkbP820ymkhe8xxI44yionfmdF74NrsJRWW9Bqxg3dLacFMU9LI7BdkNgJxgrzRPltbvdP
g2pi5Ubu7VT2G9RL0G5TADSFkbxsPzA5EIPCuCWDQqabSN5wGvILACygOav0KsxhjvdY1mN0G1rB
kEXJ+9szIzbn8A5HHNLfrNmyn0Phigsvy9n8ECeJE8a70yy3C3hpXfpjuXgfJV81+auzY9VewJ4F
wouDe4kRBjCikMSlDZmqy3jxjtveCqIrExro1mosSTzOWThJ77niBG5BUXMTmP+nQ8V/r21N7ZJz
/DKje+uZ+pftVy2sEH4bIe2eYT8MbNcTCpJfX7kuAXNPaVMzWDayZwHaAH5sSSioEAZwDwO0qiCb
wqEBKO5A8/+zjxCyJfH0MXfTvxCTdV1SwnoVVhMwixxn0PXYe2FPcORIB7K+m4LBSlVwX6PvjgQv
sY43xIUoBfPt7jpLYG+Pg9G/7r6tFC4hjIiCtCm3m/EpaQpIqll7UzwN0bj+ouN7T7YGXRuwW8cH
MMMjNGLR0ou1nhJ6LTrFXFIN6pl8owY72HaWRx0LM/RTo3V+4V2Z4pnVJQ7VMSVRYlH5XSh9wCUr
LY/5F5b8Dw17ZjP8ZDKfHRgnlJnIhyYUotrP59Lp83a683HVcMEkhtcUrykBi8GW8EEOY5B4CcrR
LT/O587uMG4weg+ggXP0ZgLN4F7exB7+9ARjLWb4HMFOOEoRuM48qs4QGtbilxFTmMODLB67l70d
rJtrokjiZmoC4WMUcmALugV2mImx/Sc8ugUJ/prmXQH4jANstyvnty4SmJpnsgBxm0GQ/DeWGQ4v
zJ8qURGbx4ROJqnxftx9XayJwq+eAUNQebeMv4Ct0a2wW/HikMIjSohAjRiEcmHwYRMqTtss9u5H
T9kNA+mPsChwxwqqrM3yt45nPEt1cB8S24bUYXo+pzkEnhqAKcrl2JF+fORtT590TMwW9yWu6iC0
q5ZemzwNAAcqUm8QTuUFCs9sTRZoTbd5jMu3XRSvm84b7h4MZ651pw/YKNDLXrrVlIGYDX6nQceP
1foc9fowAiiZ5w4ncG+HX0JwwmcFKOKv6TtorPrz3jNQLNyO2H7HHM6jTJNkBsIgjkxazj5w8OXM
WNODGYVBt1eusenPBja4wVOEtgPSC419mKZq4bkOj3IFKqZirn++/dfCTvDdNKEW6YdCFVHjoAWF
tY/mrEGLJUC8nU61iOLhPllkfzmcsU/t4qvUvvr32gKLu1Eg3xbYmNfB2WkgJ/ARU/Zxy+Cbsc2J
+Mi27TUFAmWzVrq9JvMZcmspKvDNQjVuR14mcnS0R+SsSiv+nzCfRWn23LnlWtQS2uRp/EJjjV8g
Xl4o4aczeH9CgkYDH+Fi+DXFPCeAJOpTyhHSUwuYs8FKG6MZXHPDRRRT1zoCvuUPbzeSd/Iymjjw
Ktwvg7Q2q1Qo4ZNUvSh7oNTEyi4X8hjhEbxYsKFt5jMiRS5sh9zmcwq9//ADHhl8XC5Yp+QIrMyR
c4DaEMGeD/qtrUrMa053APBc9SYUjGwLFF/ZBI2ZdF5APgJDCLQJVnsPU/0mHUm+FncqbgE//HpE
/7OCJby6OBTJh5gtbxXnP3bMUkeghbtumdOmkhalecROUFtAXIygkrD7Mc8tjBesaQRtsNQtHl3w
crFyLVbe/PCav4KJQhpaRbK9VJr6V6nsNFjFXItdypNgaEuz6iSZEXyY3BTfPC/rCHkc0fQ0WXXY
KAVdsN2owS5O1sRU+39N0vp2Jwp/1pbgfwwtzAK/wzjwjfh0onr8NTRx6LdQYnMB5rn58Vl94eNA
9zvHq9TNrdVisoZSekGNMBaZVcHbBERwQZWKAW9G2nnsdv8ePKKL9Ka1EoCh3b6yunUM2kQFT64p
h+HiduCrhXzdOHbnPH8MOIJEIESh27fGjWm9lI1mi+c2NQ7VhIZ31lmT9XkcX7iQE8EmyIqQ3DJ4
3C/3G8ugO/kBfhB926+adKM4Ub/CfkfYtapqVRqsmqhBF6ggpE2b8CqJX9tJaT/RNvJUPi7f+UD9
A+zFysjQZo72KA7KJJ06M+Rm2z2zhb6F3O5a8ZD4LtC+34kvGp8oqAFrQA/5ZUxLdqR9DVF+oTk5
D1yqymxiApa7hGQY6Hxc1XG27QeSQ5cNOTzIbIQS5C0pp4I8UcNOpfgeNYyy/1NRzlVbwXSpwOnh
caDgeE5qLweNyBRvMDtJOqNlW+FJ4TtE0kG136tqGRgPGmcyStxlVLYddlJoLPSiPwo+FgQP8f5V
S2rt8z+Wkhlz2lFXtNSNPezXOF9mwQ0MR/GWEATIoHjKgbfbo4gH+lV12Lkwyo0yWiX1bYn5WW6x
Qbfs4AZ7Y/2ZAtbjfmRFgdWRruQAvyFZg9e5h9XNxfQfacwLiJGhsQejyhQ2GZQLycihjGeoJkd5
Al8/xTVOn0FOg3Ghidiz0vqA9Rhjyv6zjanFY5f1GV1cOoeq2EVkBaGAdxCgbO9oYpACFhHrQ10I
7k42h0DPm2T51Q+pRK0tZqNE8GiTUw/90nhHF0eJOoj+I4g+J/FRlIoPacR2QYoSdtkGwaJGKh9e
QWALAGPf0EPdMIqJ8xJ+KSpWO0tVGl2/8WavHTT455PUWxa/Tvo08CrRYivME4fdZ697e4OMpMH7
8CrPMdcOKbp+9R4dsyRH9OnzIbxMJ92Cyjmd1ED0r5t12TzZtdI321xZZhEEhMiauETC6QMSjQst
N2DCHH8NFvuL/LlvqaQCHUxaLkJ50XN2Zqve02AJNHkQa9JbcJhfHj6w8nIA7QcvEOcc2nf0LZAb
cXMd+h07O3oygTv2QY351z6OMilqVee0mFCNK4z50vbEE/fVfSQRPxF5gQwnQck2piSgcM6hwjGK
Mj5xf0d2lnola+//Qyf30pRAwMNl/YMT5qEd/Uwhi+wFjRvRyb8miXA1EH0Z7yqCUmpLd91JJhx9
kfIOlj3II95G30MNE8p6uMwawvLtDTrrFMdvA0o248bci+pDrznVKHcS2feMFarlreGkLxrBqLnP
V9FF47P3fboHW4iwZxrAR17FakPm72VdXNXvU6e3ctyw7q4LnaDHBsKftNSiPXV1zPEu7ikoD+tS
YI3xVsAPr0um0V3hfiyxMd/dBm17eGVJurjYNFe034Iq5tLmdVPppknynmKYkJXFyCxMUCU1WlxO
4Ejw9NAuD/FqlFIaA7Ueifnpvq10Ny5LP9V256KjLLwykLt8nPkJ30jnaJql/ToKhlawB0lZGm69
IHakCb+uCCW8SUF8ipT0Z3WgUBMq247pYQHyX5EK6gKnxH+nL60Z8JMwlICSiCTy93CtGnTf/BLV
FGMJiGjZpjQ6OlvQoJOnRR6XFH0dp+CFyh0ZuRMzSRP6LsTa0cWAUCRzA0JaOYMfyIlUzGklJena
SdOB68XIorO93LeQvdbU8ldlneqygQjDsIXV3p1212xevcd0s0OSdPNXUms9FIkK1ZQTzSRQozUY
jmBIfjPf275FGT5vWN1N/3UpZGbPhDEYDQiSZQWpj4kEDjJ6Lv2Vy+adqQjOgpMi6SfGBMCGWyTN
DT92+cELQffQm8migT2bwXaQ7RyLU/fYOaF+hCWR10u123gRl+7ok1bBsn0qlIzigW+a5Lb75DLT
F53ccj4PuhZjQwfcxZU+buMQR2kC+Z0TReRb+a3IQsQF4ieiN9QIQiRcUeYwwMdPG6UzLLCtAqKq
NTbb+67nt8O5V4NXrkPL+qX20SNYcQlZS9CEem1J6Gb1be4TY/fKTZ48XH5rvaVljYFaxcqfZx3o
jaMbPUsw/zmGe2uxRt6U2SopNQFVB8FTWA/QK+2IGjPpmCoid2bqZORwbEviJEOnXMjguodS5oxY
uKDV1bdib/fTyI0yV5Ey1zTP9BSanNW/aJVdSgDq1DDKSKDJISgjSE6fpArSPOetYImryAnfOdha
c/AuSwwAv8s+V/2b7nWNqEMV95voQK2+g2ACLokoVtyBqMyyAYm7vvrOla4vi1A/L6XaDWMvybTh
gTWucewZHvws1TA9KfFnMKLiESuH2Hyf2RLfU3yUxnpjw56c3MUEdCyra0V1nm0aUHAFSgbtigvg
8q845LFwzFgteCN21kR2nK574qYQ0FG0UHw7XLbfU0FpOItYQMa75PsLsWslVzLk/G+iIhJ7hsCM
QZUSUoNF+dF0eDUWe5GTuC+H7xIhyxkjEjujmSHwsNnrgBM7t4ctgWWmQnDG5ZG6vqc2A+mgV+9d
rGRGaS6jLLo6Iuf7RX8LI9U6sLjm0JTX0ItwmEZglErNUs8AhGDA/vcn/STXppB/vV3DbqhDrfQL
02GQ3+f5LgoRQ+OEu2Y1sbqfMnaz51e+Dt7jFmbm2IZHerBfnJhnfZ87nIMPBSOuTMUB/VqdNwzM
HtkS37ANQPTZdXeD9ZhhwixGTFYpYwNOL6Quw8JygA2sgrOwDPHBfGGEkWHPMNWY7llUWmg+KLgu
cZYVNNNVtGsp6QjQ2uLJpBJ8CorArIPAmchhIFIn1U4XjlQM40b67uqrm4bOFAhuo7OBiGRQJT4/
nDBEhFEnykqqOPZJRbXr7/y3SRx79GZ6KYdQAB1vlW9WEVw6Pbdp4mRlwwiJn2LV/Oa/whNPIbki
PBpeWXlGgEpN6+tCaB1qjVolFC3iFru9Ih+tD5jHo72i/vtXgD+EuQq0l5aDaLxzSD1ZMDi6M0QD
SLC4gDG/DjwxoZneCcUVF76czQsWoZmZdNS6VTsoDtwG70T+ROmQUDSdGNxMwi/HxgVO+ygtE3YB
NKYf5NQePaHy0olUpLaI3roHxmy8QHb2Q6ruajJwj3gLGtR9Q0xWs5IvZuUflP6hl63xZG+BVT8A
kRa5sVs+BFwqeG2IL1ZOFD6D8ntx/CJ/4rDSTyGj8/lZa28icYSI/pAfBxkeuRu8E9A6cUTFlA9j
90DbTeeVnRvlVM478be3HoTUhwhamGl3+MLxm0Pl8+18RcpDQr7FThvFeUymLOW+qPyjsA/ZErvw
nuSJ9jObO4qTYCIk20fxF3kvjTnOgdwoRgUxpbTkkGYdV4f2n2LiBXRoo9w4O/2J7sxP9yVfRHkn
6nqsiX40OiV45aLZbSPDf8H9fpbf4rHBMrRBmSEGNknRdPyeMQquUhePb4BIy502IAlK9npafPoG
Hia+rtMASKA81aRD6CcIwW2aGnmwDNkq2Bv9AovS39mYJx0HIAkebWRRMPCwg1sKXFURuWldO253
8cXpP7JJ/BMz+famD81jm2AZCmMJRfrMNxbFZ+Yx2XKW5YWZBbMdkyPY6pK8dqhJ8bLhlbkHRo1T
f7R7NFesS9J03S3zeGhopUeed/1oI2yCT3XrWuLBbC8sblMDC8lgzv365PBDqCaSSlhanZmStd/j
fZtSZwzivl97W0QkmfKc81v3Bpj2oE+b/PyStkOGy6cE60uLHTKgNOUfFJ2pxkky6QtcZnNXaj+p
8qrslofOVprf8sfW41FyEoOQUAjTisg1KZHlQwyzk+WnnOV7jCmZQOAgqZMLnbzV3Reb8NUMzaA7
DF5yFmbzlbVqvGtDQqSnmHWIEfhUncoLJPTA27XB3TkihrTrgKYIor+NDz8lVlXE/+QX3i7iQAdp
TLWQyY9+Nyybop4UlXeelKB4Nw8obe3zBS1mnxF+mnXm0/fa71bCPd025EK8R2q6FJd1reWngv7U
gDOS0UQWPSmpi7GpXyKmgRTwt68UAUSsg9usstMiFAe4vv7AhF2YaiFh/fnoj621a5VyGH8L2+bC
n4zMFinlloc1bD4a4HbsIQ0xXFgP19HaO5BqcmINQhUPbRtkoxyNISHKt8AfXPcKAIvGveeyFhBG
IAFBV1YDba7wGqkqbewYsirXZ3FznEoDXISxyIj54Rg7G+v6HuRA5bM8G+jckrU3+Y4li2OM26fi
RkOOZLS9jPx8K1I2FsDcYe/GFLfIsahBPfAtnrk4AUl6Rz/nNDX3ryTrJXoJfHGYTf0vTjUZ9aBd
Jz95JbBVwrnv5CN5J10JBss8pPB5JvIP90VydO7w1RNtR71MUqCS33CgX1IJj9zxyAL1+jf7hKu/
mPMYEDoVyznAYPQ/N48iCa0wiSlSZGLAtPgE0nXI8BBXTmLSzSzDXW3pYR9ZmzNg4W3tmpJrnp+u
gVQdlk6iFwwe0rCk7upLiDNdBGXYWqfCLEnYdf6xWDYWXtcVLTQjaTNK5XmLpEGO/VaftnYcYd1f
iuHqGYFZ7EZWHAQ/x991jZ+cc6dfwzXPvRYUbnArMHgukjeeoosLjvLcbjJxi3fxZOgEuuT8AgGZ
AOGj2z+zISAcaF896TgG/MKQF6YcsMp3VjGtPK4sbP/3NfwQ3KHC7hra4pnXK0ANVDlLpL/arrN9
U8e8pEbHMkccop0wOQTYQPBFxAvLl79D/pYpRoLlfoxi107Znlzv119cQXY+1PXSQm76epeUC1CR
6Z43//cvvws0kI5NgKmMC45/WXmSmUE53kkzM6twmRfXzN4Syec2zzMG3YWeKB7KnCXInAA3ySbx
SgDJSJfCIZab3uRiN6dim+Xc+DWCKQ2roVdE1iTunAVTHs+wxQfXDm5m9EhnH6fGS08NCzRQSju7
4orX/sicQtykcDv8q8buKlWfczXc2WOZ4fG4ZmUEfvrolYJGBUWnF8j/xXZ0o/743VI/nZFS0rLS
J6szsYQ0A7VMBG1vkRw4ty3L6Oq5oVg9YuJI4ih9l/AAocokInb5TTX655L3SAqRf9em85Cmrzik
HScygyqTcETjTV2BAzAEQ3d/qmVKt8z/wVCcKwcHY797RPMqlYEdHdRtj/qyMp3Da1XrWMjKUdEM
UnahDtsmFSe6VxVC/sNf6WZOtL3vJXfrIsad4MczXYKn0OtCuyIjnPdO44kaDqVtcgIBH9Vnv/MA
SDsXcopBfK9jfemlMFRG5Koqt9mUH9SE0nMhS1SjDySBzJdfPXSRxdWTYzPPPZT8Ivw2H61+aVkn
0KwsXj8P1LViOxZsxs8xynOyCnrydqSXWeieu6bjnPF5gIE3TSRy9DaIA+2OA+lj/M+U8bvefKon
mqndD+koj1B2liAZHWj/yM1Hl3vsa6FS9H4vgIGkEba3+apias3Il8gAiT9QrYwW6ldRI2oAqCEk
l8ovDfBt9DYr8adrr1uJHOETYLpj9bbCFr8rrv15vTiVt8Ifxmuld3r0L41CpxjDBipL6ec5ny3V
ajj87c0vdTuYNGtVKuXhF+pzgaNZlVPLgN2G3BGTL33acBONf5qqYn8NAVdMbcBasoXzUSDskrEB
mHbrudNj9N9kAPJ39KVDylVMPkKXd4ntvA5TMhVndzGwmyk0GL1RoR6XtfYDMBbo55cgShTAMarV
NmE5mOI1kz4hqsiFd/9S1rDvqOUosrHCKV3uHY8MaJL+ruMjLRmkJhY8clzzu5VDTW4VCjrnp7OJ
0bgTXRc0H87HN9QYPpSYJgx3+g4uKPqHaAk3kmtq/R0CBMd72xZZUpazaPlYm41uN4vMeWIwxOi3
6epweauA/bnqkKj5wqqtLUvQ7rA4QqdALh73WT0ktxbfqRX4nHXyJ2yYfWjrsqzGVW1bNedWgSp2
LXJdtboYiil81Sl1e5XQT/b7Ma2ywBPBaASfRD7oTIDBei8gebwjiusm1xgBn829rEQboqnrJkCW
DIsx5FvzA8hk/StJxiiCvhTqIf1cPaiVevpaKFOyWhqhKCMZRh1hs1oJARRSI85MhISUL8M5I/BN
5mlGOk5/7FII2UQmhf7bZRXq2PWztAfIZpUZ4B7zIQL6eHtnzV69fUWzbw3B1upSVOuZNtYYq0Ul
8amQ5fAzXW1rRuj6c/RU9YqEU04KAACQ90DsE5mJj4nsZAw0XdpjCx4ozMx7YG46OyZAYRy/Bx0f
CgXv0BwanLcykKY/pisZ0MkUP9UXFUDdy65tNIAKFLJi//+N5MQBn0W5D13a/UC9Bn+ge5NQiOq0
vHxgR21Uu11kHZpNuh//u0QRLy3RFm0sHGkCM2cHKO9ZzDSAdqXX1Wrf6YNnNl9u6U/riPUoN0Tl
sjfx9kAoU8yqoXMlmzES+wusDGGMpHlupDuWBaaHwuqhvQE0Yx2d1RkyHpVvFRcSTD08Q6uJ+F+u
1znGmypa+HQEj9zhiNCspXg7ikHxeO+HZcyzhK5G1B5n+6XWaverDmPMwX719d7nTdEePkWopnPN
izljCSWHg1Ak5Sd3UBHowj4U4+0ZO7LR/Ta7bTl3cElFzqI3+YF219xz2F2++elZlMSbk3j9StKo
TUi8DjXtvy0u/auO/rk/s/b86TfWaFt8RPgWr5RCr0Dipoak9/lpK5OrD1BNucK1RTaxYgtdlXJC
liNETryjI1gz0Wbg72dp/C5X0xK7q4lE4x+EVWoqcVLzqGngna6jvUTRLFwVW4FwRfeD0aSNgg4L
exRQBrpqDYMzMxXlCARKGKUt7DmU1Cc7bZA3uHPCchIQf/xAmhipFRODli742AsCUYV/WsDjXx1j
id8Qm6r3QaMEjdZPXkDaDONHi2ykWcAlStEDKbGCI89nY/fSCLDbJ7pMHu2NL5QH9b5qsCyr5Cpy
AlsyW69oMyuL50ODOz+wBBEl4Aa3uDYLj/ggzsZfVKc9U4bnjIyzOeuX6TvFN5OdP7BRQYvZs4Tg
Dq8DKBQnxpzMEvWzidskI2+ClVNImOyYE/e5ZU3vggQDA/ivjUBphAkJE+wMFyhFRxCy5/nghFiN
V8CztuHa3UZZxxrQLcDrxyIZlLFfpX7U0MPaKzlDDLQlO0aPvVVa6lbjI3umAxyiweqLMBsIXSIW
FHNXMroyi4UZONUbCpSBqN87ZNFqYcHp1OFKHaMDAvyC9biJ+7QtY4aTZCLzPgORny+mCLCVpWLr
49G/E70MBfoicEU6/Ege/D1mkusuWolG5V52eGiwJaPu4LQItw6WccQxivbxADSVsoAt5cJTZCHI
zp+tgsFuK1PGOrinBBM2GBAenmq/Lh1BDfGcpLZtUuTsFnTkESf70w45TWsvsmMsQiTafApldN6H
4OXfOoQ2ohgYntazutUhTR9vpAVr2IycBsqmowJBDrq1oraI+5dDJAXfTvvvXjPOm/o2hX/6r94P
rTAvwSu1UGVXzCOZiIakAf0Hs+5UvRDDBKDwLzX5nCC2xhD0itNm/FTt1PieOqWcy1jkYugq0VUp
9oZhQkA0jjl2Hm6GSxiz3Bg3GlsjsGpPUA0dTXPVLipbdSWqwN1oyxyhXzRV7xz81s09SWiz+nEW
1EC3tfyTNs6bqO8skxt5VHsvVthVhdP0TDhodZMnMu3Lqee7PVcIIxG9W6vbxRzcdW18kQekR5rg
o0haOGDPAEkAAZogAWDSBvKKTxIIttB+zzII0grDbaVCYRsr2qmDUK04EySdT1bF3BxE+aFozRp+
wqqRMiS57adgZUx1kWHN0AVCrFaOgfJUtqspGmCS5focFNXqpkrThSzopN8Z3oNHt8UPjESiZZlG
Es7yugdUtW9UsESh8N1o+Eh0fg5SrmCCnj+yCfoVcV2h2LFoDY8agj/fNsARxDTjpHXXXEabCqLf
rK57wpRCWGDcGhjsOYrGXWweTRTZZoO33syVEVoiRD3UXYvLoC2nNHno+wZ2mrN2dohBlmh86W7x
5Ynl+O7wXdX5CvAAgxy5mZ+3/WC/CYzxpEHHTm6ivK7auCEsPvtpNcjoH8E1P21UXrR9GwX2olhw
xYevYu3TlauCpuyca8CxEJ6balQqsBLNjgYvSE8Ga3JJADhk4c9Xf0nTenS5zV3FkXcK3ejXxwyi
OIGRV5NJJqAHGpVYTVgAlHWQU/pmRocKjJ3WzPlBnKYydAXNl4n0Wfu1SvlHdvKc/IvAf5xkHeHe
DgxT7t1BRogRpJpej8hqFhF+wfRQ/mAa7REul0uhux98QP13qPcwNAwTBB7oz8/5jyPZZZzemlsp
BiHUYWJD1FjcRNk4bYp5f4Ay7B67LTZ/HZvnl/AIsAfLNaK521lFbvginA4v/PBscbFr+JDlKFT/
GlSK+L3HplLlVl8MWmORgao8ZSmKg19SWSfyr02Ks44phKs44g/iRUIvG0JJzWkhTTm2tIg5l6cK
NuDma8q/5FletpOz5bWccZybvJmaP4ddhA7N4NZH9s6K5wbcFSVwIsylvsDl7T3UCCZSgKcBU/nZ
8Fc+M+5a9EmWVKTVT3FNdBGiwUKIs0tk3Tnv5YKAzBXbLyMdMCxJ2hcn5CMfAGKn0BPi1zKk6jb3
Z+BK+t0LbaPF1BZk/FFbYQxeFa1crZqr62d0VhRABTAhxbg2UlhFOBt0HQ1revlghNRHd7tkeMSD
UxKDqsqpzV2gtlyIQgRl/VSYB9l7jCn1KYHD1UGk0io+rVq43fC7Qbss7KWYEZBjnjr0CE/YFmNg
xytcgmxyQH6kNP9J9E5BHbPHp9ymAA7vW14lQ9vqW/6kFPwhlRyieYeLOnW/qEZfBjyW3l5di9dR
mReZ8m/s12uTWXiXRRRBS2X+tCiW8G5g2Ysc4Trb4uzmtHZVgBKRYNgkEpzTzEKwl798e/w11ZGV
1iFNwX0zG6Sbl1hgP1uvErrF8G6jyLBULv5pE1iiyXwM0rP5iNywifqAN2lYwEu6B1LHa3BQ5hjY
VQfvbfhUv77VdC6IHL3o0azPEjZHhEriOnW2GCSBhfDTRm04yZwp0I4YGlw0dYL5Txqg6+FWDvT6
F+PsfRTM8C1G+5ylWzJFoFgusUzX+1Y/YYqOcFI22LbUVARoa5ELI90Jg+FPXfEDSy6MV8UUmRo/
KAWW/jmvk+rBTQMfFzZsk+x0VghXENO9qa8ZVXIPzCRL+Sw6KLsQttuia+zuDZOmFG2hwEZj02AZ
mf1OUfnwbqX1xLAEecTTj8gK3zO+g7AoNM2aIO2MUHTjXxBacglm/oMTlx/rgt5B7vWVPsQQeDCD
pgznODEGiQr3gOF7jJH47Dk0zbH984ONzu6Cz6Gx+EX6upx8bW34rvE1hyUsgqZTX9yCwVScBVZ7
JV/ioi6sQ4d7kbG6b8Rx1G1RUoDZwoi1ZJC574Y++77nxrvnzcXZPwCIVvksjGZ2v1zq5WjYY6ym
snE0iUMW7YGf83IH5fNhcecd2Itx8Mi8Zo4f9bDjWs4qKxsO/xf/l1Riow6fiYkulmnxoEWDjRoB
XeAC5QFbpmH5UiMFICHsD0TZnxLh9rONaC2sx5xfJE+UXEQvaQNXy9ygaNg1RKv7AN933P5km6GH
UyKPOOVtGm+CBHvmW8E9+GzXJXW8mmr9EenbeCeHj5GDz+kDrgtwzA8EO6DaW/Shpyd5tExaeAC5
KNqsRFcyVkSzDvJjbFBaWnqj673VdfnTbs06sku7LTq5s3Ahj4FK/XDo6CEnt33oPTbLM6GZWiRL
R9Z0DvojuLwKt6XSv04DmxTOLA6jMJ/JgRfrmThxu6Y3CyGn92/j5ZPNtqgA/1ZFdVtGPnSDYgiy
85XD3fdjoAkQy7jdsw2Emdr9kDHkni9jHMkP6Pm6fYHjnhUoNUoxnxt3RsbGVmKS3Rb0X+zBxXUm
1i3LUmp3Thwh2HjVct2LsnloJlhMjdrJeL5J3jH4e21OtrvCvg7cOHwD/nDEcbvRjPf3p7osR9U0
pMowY0gJX02tLWg5f5wQGsDCOA9VcFkcQhuz3VOb/nXX5+kiaUBFMNtHH4cIPdz/hwrmqNn/8P5Z
Ng47khyGP/+TC+gm6z9CxsPXmY0Jmf10fqO4mSVwBSPhJVpv/nBSCaoxM7mUKFesGNqXYEZHeaoK
ZlK2UwMyb5un+sPIr5W1Iu5utM1QjFNbpm9YqCFXt7OfbFYRy4XGqkgVaIhQ1IcCZXaoEue4Vzz+
3F7SCuucw6rLajAWoPbXSEI8kjjvi/k8TAmGR77JJgPbDBWU8maHy7zXA/4drOiyuVkYI5du+ZYF
aCzVJE+CZTXn9kbkh8iKuCeiHHZEtlplQ4MJGZDAg+Z8d4IIH5kQYc2gbeM/A63s1JFWaZjoj/px
cjsGfBSDJbbbe425ekfLzCmJdpNEfPntRqZrOHvFurFrC9Gxq5EqCCphKTPuqKUgpVNfZjF7v4yy
Jj2KKBgUqjimazb7S9GsKK7iprTHwc5NjNAsC6lLhR6LDidZVN+V/25JYlg5Vw9+PX0lxU8saxTR
FQVRakY+KnFNWd+/8YsNv+lT5BuMEcl3OGdFP3GTRCARkvYwMLP94yr9/Vfo/6QCrYBnZ9Al+wsB
SBiq5DhKKHW+omq8AtAg2SVRqpsU6P/M34Rjqj9CPGdJtcKb7yI7pIba0Cy+yAIruxLtMbnTkC0E
pp/2+5wykaTgJ2ar1aBH+blpyB/tQzV/EO8uqQNfz9ZGlGdLA5mHHDV94YegQZhiGiSgz4lGOU0+
pc86BGG0Fg+qNKdC+v4TmD59uQ4Y2hFecLZ1Kc9GCEUo3sXWCdOf8vsJws4834QLqIcEhSlk0z4+
Fz2D4bISxxH982EiIA4ILXSmYS0YEUJZuMqOywZf1cbgXugWCu0kt+kTquT9Fml0s7YlTWuFdLXx
m8Hh7/oh+L8qL4EESCiACWlbLcZVNqhzrrlPzmQmopZrXnJKn08Gr76eNosxlb2s/5MKVs+ILtG4
MKzRqpd+cb8hyE2U9aJnQEqGblEV0WiNZ/qg5+b0rN3USxTUy7bBfPG+f8BfELjRXnNGgQ0R5EQB
J+cVb+V0vbH9B/fOhKq5rNEkhw2ELfZ2/9VY/Kg641Es/9nFz6Mqnm3wLsGSHd8zEZMqBavLaPeG
x7N2l+gOIcU1V+34kVQV4tCLWdvVLBRcZhvzoDd30DaqH42qOER8mF/b2Z5Hxjs4jlXj2Banr0Bh
ObCDUVlL6xuo9uhhr7d6UfDZ6EzhXZ/lHxVkn4VN81WMO22aSl6VQd1bgOFQZx3AScmh93u5w3gQ
5VCUyTz4sfRq6r2mO0u+fs2wGHAzjT6s166TZtKsXI/2Cw9twpW4YaGKWYEe2tMly+lpAmAgvrZE
UolxszLCArgHyK+DXKQN4lRKU7KByEog8fs0sQm3U2zGMZVF7ecOlFL8ElwF+cYi3Obi6FyJZ3CF
98hIG9Mi4NUJh+Kl8ALPiDnVFo2dL5nJANNW7yWhLfiP5Go3gpFtG/J9g1ghP/afoRaX5lpHOOOO
7uXnXOIC+6CGIm6dE7a6ciP/9tu8/k+Ou8EVGb1iyVGJTYUWd267M88gvxPaglpv9VBcLG6w8Wb5
JcNL3sQ93ryRuWf+Flg6hrDmcL0ZaZKbhM2d6KSW/1uNvH6FjkmCE1ZzXAWhmBitFlNIlynjxgDx
eATjo3J+/BosdpzMNfw1UvssU+1vhVISQxGRynYYggl5Ge5sK6kWf+TL5yLnJ4bL5/sdEKg8WVW8
4FmKJVpCO6kBMiAm7rW55UNByzJKL2OMRpBIwho4yePF/7BExRMI2lZquF/H9Zd5v4W+q6WyQlO0
LtBJj3ifb/DNOunuP2yf3K2T8D6lI2diBZz54D622rcUtLnMlfCZ783RvMXH2HJ5klo3tlMISUNN
zs9GeNW1pa/tOohnAdGZsKvUo6MrEaZPRTcQHXoOSJwM+wQxKvcUjxR9XMk+WQ7d6+5Ex3NzFdW2
iFtosFKReRbLrt5x4+MaR70CBP6aBnT+81wTiULJolv3roaMHxK0Ed8msr8pw3gK88KqIuQAZO1m
W0UhD4cBwTnwha+aG5mWN6EIQwqWx/CztzgDjs+m85/+N+BJd5mX54wfcix3oMffByfZH5wgXXf6
nS9sjcUuMcjHksKmDREGbqb3wZ4+8124HREElDnyjOc+CoIKLlxWfTctgGAgEIbH2kRVbU0g3NHD
rpNUQG9HuuC6IDcz4nU/zz/0A69A5nc0CTC0ap/Op2EBUekwe1gJt9ytMAoGZHlEk6sH2UneGYuh
9eR8CRLQreOT4UTTGf+KDqmfx3JhWRcFKwNGvn6bzLDA1SXTmmZylp6EqhGZnTrC0rscN1FLOZRH
6RA3DaEThKlv4IpeicpUKh88DEzKXfqyFMAeq5sBUHiUSfP1PGH95I1cVn1flKDF96KOWz45Zi8M
J1pT3SbeV939V7s/bNnURkUvBkmCMkIR6MjFnTL0QOot4W0GfNo6xHD03Lq1cU88EB6KGh3RQXB8
3oyWUnt+Iy0efOGiJxwHRHc+sretSapFFDPFOM0gYTkJqU11EMuY5+qZdQRiHnIHmVSDsHMEBrkX
AixgibWITspEhsvu/R9aN0ak6L7cIkY7BL0L25EyHu5OsVuYjftRtiiVR6JaKgTRtwQL+PcrB7C3
/Lus7yoAQmaGA2hR9vD3jLyeL7XPAqzUxPT9YfbQXV2Y3WTrf2fndE/Kg6N5Vvz53fqPdqRAuLYP
tnoDeSZiwIFQRP/RSABFuc8K2gNap/gG1mA9SzNHS5NIlFQA3jf8yBJG80q7SP24ZQC3I2LHnHjt
jW7IwWxX7AS4/P1d4+qGgNhgb2U2vOifCPw9Ej+y7IfV9a8w4mV1phBKMElwMVhH++M78oQu8RZz
wqU0Bk9WC8HoMZRZte2wLkMyHmzPeT7TzNK+0fmfEDyAOQIvqCeMmgBzf3LsbibjJx02Lxg8316Y
3yPBxNanrBorumGZACaRlHG+iOoluDAFsuF2YTM8zYHxuB3gDg+z5SiePVc8V9Pzr9DBVmz6ZM+2
496pRqcDJd19edMxbXq3pPXyTggNIzjIFYOeAuKmJfsHP5WX5PnsEaAuqpiB0vcHrs4ScfbO+FCs
d5FnHR30MHXRqxVLUr4w6qEoTi+bYa1GaSXL17VgiBhC0gA5NmRQpgw9Z404eKL/BtJW81ohfwRN
gm9aeOMV6NcDIF6o/7tX3xiOw9xTm0/yPzXuoT8UBVerDvLWa6PlWSst47kA9FXqtprs7Jg+xKCa
2KFV1ST9bZUEBJokpfM4TBFBM02wkglao5T15VPIqLjG4dCng4KNRtFvFcu7Pw+nNzUelKbGI8h6
EdR6O3K06SfBF40+265f2SuxeJ0FGZPZThOiJpd0ZSNqwd3VnCmhm1RkG44foKwHtAfnnst6TeFJ
LGkuA5hU6ydsY6jYMQlcc5x0l8RsdcxJsUbxOnEHqdRMipI+ojhU4+JIxw2DZdDhUrQveDUFOaCc
xKrFIsYXiz/nL+QaZxhe8YI9lryxOhTyZpGAIx2d9U0+kUUIp42JZB47dtMUstQCLC0x/UrOU7+U
qY9OJIdpfdHWzE6jnKzfLq/4ujuwamCAnXBW7TZYN+tjT1DFVRGxTRQLfydG+19iN/HzAzSlWl8n
ZkiFvACLplPlGdbAsth3hFMYDGrpijJfc2Po5uE1retCMOPHMzpCiy035MOV7k5Xv28PSfMu2R+9
Z0kNZC/jksGC3mWF3jeiOhVX6YJNaPW4295ekeLofzoMRM24cZJ3tpS9LCYyNDXXZnWncFmvSe5Y
lbtXR5qpsUwssgKKrIh2fjq/3ULkJJGAbNwXIovI2f3d36jVHK1qc3GOb7ZT5UODm1htQfrbuppy
zMOOqtfltuUB82W9UPNulwr3S5/ap11rFprVSknjVjAKu12yLwrG0bKsiRn8XWMMQedsgulaaDvk
aANK7g6FYewsEaPkL0BdOHkZ8fiCcTW4P1kDcEZqI7yyTirgeREO4d9MSugjY8KY4gL6rklmYzw+
WggtQW+uXeme9aKfo8CDOL4/HixgGS64ZqeWm30yXiB1lnGmjd+9XjnFmWiQG9cF4hiBSwLag4Fh
3i687I2hoUzI1xWPnoMroB3KV/OrAqOI9HI0ueoSnxrjlNERyvPGNYlHZNpLqt5vfVq/E26Z9iKn
R4o9EIbn7WfbInKIFjLbJ0+eI7+ZS6HW22VrRycR/r+CYHS/VVmHVItGzUCL4q0kvVo7kcrtvORs
Awz3Qyz/kuTWOTh31r6nn9rHcb57ilw1ftDdt+5i/lIVcx6I1M8h9/nFjdRzQ2gRGLVq1t3HKHTW
kT0pp4Fq6cmsgIydi+DH498tu5oUxCSbWYHP0iwSckK3rIMJVxcJFa+awbSoQW4eVcPf9plBAP9M
4y2Uhfjo3EcgnrRbgCkE5PmDTMLqBgcryLt9GTFsdN12e02qq1ikA1990oVE6p085ypFqQFWVweu
e7BhfxWPEDBb5qi/eM2WlBWiViXCZBuYkk4jf3HTvyDGSirLEuDiAKrG7PVpRoULObMNM7mDxhG7
Vdfn8A6Gyh221+aL9Cd1TNRGdx5RQanjzcv9Kmw8GduChYhyCaLBPI9RTq/qIbhjnSIq109y69Wn
0HFpHGhf3fRqENmQjOcCvejpTDLaGZBtBISLgQ7XNA9TgG9w6HGMKUthCQfzRiwz7aIH66WGVb35
oCLv/SooQgef5av75H908L53MHgORd7B5E/hX+EppMHXa3FTFBgQrUKfg5EiPJk73N72ptULa8Pw
MbdOuQiLlU+i8+jDxAuOhww87j654aNrbgMJnPaUZMs+kYB6Y8+M0GWEn2jLZKfFAtQxZ6/3lO60
fXz2mBxI7/1xqdKgrCgGzzDgUAhBEHCgqWkPrjaY43f1Jvxh58HSiADsVKlXqG2kOdDRKVckl3GQ
oIdVmasWMGTFtuUEA8l38RObVJOXgYiqfHdqrSXulR5IYrIkM91Kkec8yelXBac0DWZA9F6PRGQ4
6GltPtJa9BmrzxWD+TnlVR9hzYUhU/xt6r+fIhLe/ALdAR7ClCw1NTzRzU6eAuaPSaLGgTfn7ZFp
qtu/j3Vj2Lhdu/+KgQnBy9R7scA16QDA1FtpJK0fMCPLATXnLOiFvk5vtLnxfvlkNCrRVQThrIxw
R88FZsLw0aYXP4VswfF8bDJMj/JoWvTagYHnleByuvjI7jyzhk6coeyD569GB57L9qfNaQOaMVPh
3DQngpRN57h/qGzpLnA0AQLBFMHz9GNKhLwKKdaa8OhpgjQ9os0CXUxhangj+rwoElKhsJbAe9he
AAPg+/SPslfiHD3fhDRv+Q+2wv5K60IKLWd6MWyGWC0qkIp8o5FoOPcrCmgeAD32gvvqypMqhFv9
wa03Q+VIjcZuH9Wx/L/1rBrdNBWQTHNnmHBtwGb4Ftzmlst/RCyH7rwDFt74dWTMJcIcfUOix+Wj
d2DVY6/ZDKDO8w8CqF13zNzkjBv2XgW+qT4zj2MRoQAXbII4cp1zCboUnTLFu6vmJadqYtlkvsxv
f3HmJ7UY14JR0fZEc0KJUkmd3FjoRj25Wzsm+7qu1LtzRyqnnECP3Il82WVG++QrsYfUo00ISyw7
iNUXsorM5tazoJiwl8hQyI4JBsdK3DO08OsPNDlqdeCu5UTwN2n0p1XbE1palbodu+WoT5vzjkTk
ZDwluzUZnElwWclJCge134FpAOrkyrL/DTyjJOaGp/uKXGdkU3Maztxd2gG0KTZkk/c7VLd5IwRC
VbNvTzpE9C3N2u071D5dvT0bwAFwfRRJaU8EQj+84f+MjnKWs7BvTFef2Ci3Gzj1zy37/oDGg0ns
I9DUyRYVbammTYXianATtr2k44Yq/H2mrZhEXQlN0uzpltV8hMGKWibjiHmDiNfLs7oCqs4oietN
cPxRmXmEfignvly7l4MMV4rTmmJtLQeQs1ZVbiyytVUBIrhBkLcf07GsBwcz+Z3xFEIhbp5ZCMK3
cXQfgErXnSgU7+jZUPQb64USOAPrhUzsnqfh3TT3C41yLpLfcIXWFW284jgf/nE/OrRZb1NlxDsv
jm9upbshLoWjavm+4rnPoaXxHJ0NHE7/AduwneQlUzFLREwhn6r+8Ni2WS7aM+bIMUUaeh/NfW7r
OB4dQiL4neYcLXQ/xDKhadMdqX9A+9fDvNME27D16G49VbLvZX1iyRJoRtpQHhdgvlj99jEOyHx8
2IpUtcIrWEDiqcDD0ID1IdoLPT9nvjY/Ve9v2XCE3gmmWpP/piX1UqWLDFABoUafjG7EkpNcPJfF
N7YCESkRDI+SLDmtsSxJ90kCNUt2I1M2JOWBCxUz+qaCiCuB0LhK4eH8s+okgtMCB7cLG+hK69zr
6X7Ft7yPysUVEm2n++vHPPNkjYJyNjcGRfI4a3dQoN6GkTPXTpcSItRVeXg7iHQLmpQzvtQflziT
iJrB0nuyJniFN4jY7Cu7GMP2rCcjsScxx4Ap0Tw0hCwqB75OmB4kFlO/3ibViI2phfJN4StypPcJ
XbGPyPiFq0ND43l09RmJJ5UrGdUBU+ww0s5LGZfzA/wsVS1Px2sI1GYi1QrWvpTQBlq+PE4yAUZr
n2m8HgDLrkzjPZDIicJ0rfWuq+lTcr2F1V7PDqr6BemxG4CB1Y8MSp2aRmpD2taxxPov/090HqG/
IJvK/fjPMrM4Ltyf2LYM6/Unat+QHtmFXmnvf2uULqflG558PdDkHNrBuyywCfltEj2vuOahr8Iz
MDepOQNSuLLRlnvuMoasq6BKp/QtsTPQh408yoiiF+PNxw5PVvzPDIsDG/5KgdvFbM29+d4/NQ9E
M7h3ireCPet/5YPsZ1JemFOckFewJ0UaB7+AkjdTk7VGF3Gn7mcYY80DDZto/ophrg6uqnN3usp4
W8gUdKPaI6531IPAhb29/Lv+q/hxePNHPCZjIdR9WxF/ePUHx6xuLGgN+tg8GqjMMS/ujed3RR8d
me/0vMeMeZlvidhCVwRP0MaSvfh4tMHJg8Z2R14BokwaKxVqpNn2f2ci0GBjEOmykMNG4gUZqc1k
dw3qKKSdYqMJCyuXG4FTeokbSp4ev3YwYrAlfwBTkNliC1iiV1WSKdjLun+rzJZgxwLbv5Tf+S27
rEGyKHuCLoLQ9azB1mSgSevdoglMLlHbuehpsc/D1XijWYti2+DtXKEKLdbQvNSGtIQGOzUXnskL
cTxkoebwaJADMO+bFDjYgJPYaVbsKDty17PeOKOj6zL6UL//U12h6IsKPND5vXHocHqV0XfcmjSj
nxbJeFqgOJuT0sgDsf/ar9ktaphiEyAahRRClynayGlw6xT3BBazSNJ8hoyDkNCHoglrVy8JIXmd
coPiT3VmBIsnuHTJ1zU/gz2FO7j3Qv9XXrGpzn848hjhwXUkR0iOeNstN7ZWvSeUd+OGJDwQ1PZB
+LWUb0befhEcmzXH87T4uXODPorVF9ODQln1GD5ZSqBE1E6H7qJkAx0YrXq+g4XZnv9TjGle9a8o
cWgk79azMW2JIq6spzzkEqOPs9NWB+cp1PDurF712FSflcTS1HBCdBcOP0zQlBRLHt/D24K53DVM
mavvLx6yHlTkt7fEsi+HWRiq0F7WIxJjOeNorqUMUG/D4eEuIgBejslur6GzIXyeQzBZnMCUVP8u
rD9mVbf7vgMMyvnyVLoqR3LGqejR9KFEpnAKVzrMu5gF0X9RBE2Ui22JYR3NIjgpKgUm3fGw25cz
ytwJr3l9UWGXCU+Hvrp4uO+Vdb2ck7FEsYjwi+/YZ7iUtZ9D9FkMN1S2WMO1OuA3HugWgYa5suw2
WfHsDS9uzlNmJ/ddQ16DQ91W93A/3NceJ6jeid9wmdn4b3qxZgOTxCUO5dQsv1DqLcoEpe14dG6L
IFKDJcSyIgrT780daEdKEMNRp9qOA/0kPnqpsdiTZSpqq5p2SHRnHeCZWnS/UROmENHNW+6GyKpN
Jwa6xPCcMMmQcViYa98T09VlfVU6fixqgxoBQ7cQB5VmDG4KlYInSW2gC3ii5L6oy6bPXivphDOI
fL2l0kBA1blCOdoZcasASt9E6/b7YOgSw3OqTtrCesmxD4QuQLGywd32wRO8L4eKzx0vOv7df/xM
9c+a2KtlBnpn5zMafFBjN465Ren1TIinLyTQdruQpm+ApojR6cJBsED3z6d2Y7YqhBki3cjDc1re
8jirbKVXDvgaFVnScEsDpYNVg3DeGPeCadXp0UdzIA0blvcAUDoHthw+8qwp+udFxRNk0qhwdnem
uW2m9sfzkGtl2pKo6BMGkg/vSjlkspeG3/vn++KzruIp2iqSpAAMIU0jSpa5G6fdnwoDZ+tpWW2f
uAjOKIGj2qE1tKnjGJBDUhvJ9349MClYBQpSgmWSu6W3e36PkW3j0hgzbmVsxf+OSYhrEXPdb99z
UUUlxR8jYqcdYkmsy5DbYioSB5nrUDoRpmFfAYYsB7qjUkn4b+8JQ55l3EolX4J2n1Is01rvTaH6
SeKvUpMvBEInk/2GQ51KvjceWXe6l7qNCUkg8Kr7s7LVioDXxv3ogIiFvgAcnWI3AvrPzduFApxQ
0pZbT1Dy5gyup4TlpibW5zqXd+bEJmj20wCbWvs9TmLrQhimZQkTnrEXxYrbaqfxfj1H+bkF9GI/
u89AeQzKaud5JgRpff92QRINmanexQvJM4XG9C3OhE2N8B8je5SakMvh7Nc7acJM7BSv8Zc/UBy/
5nydFJBb512+YNDNwrHl1qC5DvM37NBDMFyCJd0PsQOpHHWYsp9Zc+xrJm7RRtnaHzohUBA7JSRT
qQKG2lbbAmb5Q+chfUSDkXoBSgCx1dDKDKzipuIQ890N8VViGJBXtdEvCdwvuQ5Xj3zHD/4ZJbEG
sxcDQY55uuqEMY9rsHkM5PvYnBynQVc4wWkL/FWwAhmtsb52fzaJO8cVjAzHq31SpUboQYJcA6gA
zIe2hwt5r19tEAn+kbsoiihcun0rA70EzeNkdx0yq/HHO25j0UICfpdotkzCupl8IU20lcqMjw+U
tShkpxYXtNAMV7QcT9gxAjR0iUdlTDtfKBUMNc57diWNVFPIVmJL/V4hbZpxfH3zwRD6/mhl9pWI
eEumEZlemUOqrjFHtZxpOIfjoYbKbd/JSkSOdfHkNPyRFFdZCNjtcSv1bEOSlMUiB07jjfNnt8/T
fmLsg4sbft+1Bw/0oPvk6IGpbyun9XGhc8iE9qyN9aHEldN7PKZvm6jDoTp9BZsYEwd1q0tbpKdn
vCUen/k2Tazdi++ObVuFJ72DDFezU/TTNJnEZcHBbBBUh/ywme4busxpz7HUs3OyaAtx8ew1ZUeC
Z+8VBE1yBhCDenq0fEgzqmklVam0Gegt6Iomfae/AIgyAMV/LqY9wic6bq7FI0UnB8QQxA9kY8mt
ZeODkXt0fbk6G/uIVm4FlzJvaVbAt3g0iR8UFrqgln9Y0JEi/mDljSrBP5I6vMbO7/4l+DDd9BaU
F8jcqLAAcG8mbuGs9OE0gvNtbIeoCcBcCDx/Hs1Wn/QwuMVhI/qHXGsGYFUTVz+q/9uTRVr7c7ii
Cg9v0IhraEVuFjstJam0Hs5/GJGeESNaWy13XaKwJ7cFhWWC08giTm3OrGjjtu9YpfwpdVGBYnYG
xH4v0pJExoJBvFdjkOfhqEsITbo9l7QjkWkLQZBYOs6WJb5+Bc8atBKq/stgDnLXOz7prkvrIGyl
sDW6guyQMyl6LVaWdazo14mzsS2XKVxeHe2gvGJgfwk8b/Yk3o1lrMNrg4Cfcu+n/msi1K898Amb
EH0wpr++YVjWnhygDA8CMb/spdtcp86RDNpEYO7VEdywoWjeBtBgrksVwwdPBexCd3jmPMRQZ+ce
GTshyxKaEMl3qeHot2+2bCht6u9XsjPumKdyAVUS/dpSTCgb2P7+EXjy32LcxfYELc1t3S+DK698
9LNs04kcndiYsAl+SrVRsG9s/tt0pD7JCbN42cUYzFDTzaG1ZVAuMkqpQ+6NjAI5zyVQj8qVzV1q
TGdD0/jOiCO0qeHtXnw6H8r6oYTnRC8KlkwMaDYlmeqdYRYQCOGyu3Q9HQjnfx/QhGVeXqJC1Eyf
SQ89br6Cs8x0AKLOUiPgJKAkFDEAlriUIWj/JPQJVaFKJPgh29NMFnyoWDzGn49CJaPgEKpO4jF3
6BOfJUn867k3uz43/v4Ys48iTap0XiqjzD0V4fteskVc02iEKrHvTXKK/4ZLrVJRzgijYmYMBMuR
qhNKT6KWyyJ+4pcVNRmGe5FtYQCJ+G2vWUx4kD1WX4I6fLwuEBLJZjB/mfMaD7apWacd4qhnjIk+
z1W/8Sw3SlnHFl1hxZ8gJI4Y7yckF5psiGYB/fbulyKN5h/2kUvd/kItvUc4sIR0bLUGzdMSb57n
aAgeq8vdSIzuZnyXBYfsSi7wyVRi5+Yu09ise22PjzcVlGL0Fvdt+F9mwSyi3knksO8Up4bvGFpx
bfqJrXxNt6i9l70pEpe9itIvS8rZCrtfI9pBopFWSVQLPyC7m/irmCKHH2lu8LMg0quk8c1iddEY
stFn8TVeo/iDJrpwZhbbNbE8SJYYjwA00HmuLxSKeJYaUQAZXub+fkhDoLrSLfxZ376v6tBw2bcq
WG1y8QMe4DLjjfHyBWTIpQ5MTX10vkQc1ReIMKjGgfYbRt3Mb6WJnKap76a/tmMmcVFo47hvklWv
TLG9n4d/+ELa3z+/0RXO0ahdsqF08W78dFU917oRYmNhjbfQzfx1jhhJEeT96wEn6aF78t6dViPA
+EY4AeGUk8amPMTV695pNrFJoE7j5tJEXTzA4Hi2uSnjZHGT9iVoM/LwgJjnLnDrtTvnStjNM8rO
zLd4qyrnBUaPJwDUGjvE0FdVTzB2TrmwcQdJdzlObjFDOVv569QV06eDzT0D6+kvZWYmt7Pliqxk
Xd3rrOwugkO5eiC/WXD6aTzLfu5ZVMfIlTnekLC9TVcs7w8OwucUHwwDf9fmNYqHfpwL/LUKRDG/
8PJmkGgHomFeKFUEkhKHirEsnEY+meEE3/94wP8gJ2s6h+xQONzMuvxGz9ed8rTPFteezESQ5jzA
VFex+4iguD+9J3/FCdi6RHzpZcYSoKr+O5BHpqKSvITLmNprQ1hFdTdegcl74XGAU/b4eXo6NvgY
PC37pZsNUOVnmx/OFRcg7quaKwUVApGCneFoN7FS/zWrrsBWMEy+zGcMbqLlQpI5jWa9OiEwk4Sv
XdtrR0qkUdRuF15GJ1a6NOIM301mbRM1HSS0Sw9L4ZQrHlToxQisLfIwgPx2rmqZ6DB5FEgjC7yX
bRNGaQ7dth/nD7q/cwtJH0JKshtSskaArZ8Rirv2x8M8NSKdCbFDr/ABqMWpyNbn+yWhRfJBV3rX
Xegx/eRTSNfvqE2ljRsLV5nwHhirHelqPOjN8DAdLGdXrTXlY2VPWN6EtSDwYUpBKYx6aPcPWSiG
Pt3BRJm9hT5uQZBqW0bw4q90YTYLJQPE6OaU5X1ht4UTE/FgDPQhEKaKqLy6wwF1JylKU6gj7Tm6
AgcxS4CU+eISBScRzLLK0diNOrmZIXL5rU0Fl0DLr2KJVyryXPM2KVQYdIKvqPt7bCb8IHVgNR15
Z/opMJ/WH2issC1psKs5NennhQaj0pNxhS0AMRuYopxm+iRMkhBeKSLhiF8BqqOFm8PGSo+Mb93z
hK2l4012mMrRoj8st7Luf6zaa3KhkSO7++kpilyuTmRHcckKjz9Wsg11pgxTbZSlcOUp8uc6ubwK
O6jZSP97FmQcYRNiuFZ4Q7WF0ISkXZyEE/PCK0n+fIX/1dX4xRIV5UltpWvhwuYpUjl9T6fxF2hF
CnnbeYCblsBaq7kAQOpu85yogU/DzXgx7Yf5OiDM55EWFz8XQkKhj9svAuWoOhp6vfhz5Vz/Zpk3
sYMF0RRO52ssvpH6EuPQNsQAHPqHMGeTTdHORmxHYTJUQDQ+yg1gD5Y244Lm0wfwqfcQSc43LjQ5
hveHs+feuaoQr3PmhO4ktWE0qlk1OGh0v03nQ2K7HhwIE6yx3IYW9yn0NLOTGx9iO8kCKKkaISh5
qzOWbNHmM66QDJmoyAXtV26+R74vhHKVdrR4XBPxhJ3CD6mCdqzWu5xNm17PgyR05K19EUvr0/n5
l2aOFpYCm1IvetqD3I90OYsKpdfTjj6/8w4TeWEwg3CSeLCnLr4tVAzQSPO6h3SpK9eE0HDe13Az
m+MEUgkUoFZFslspkdpL9Ne9gPlKL1hrGYqjLvECJG3/LkHjjywVJabXB5G6/HQxKq5PUNsms2qZ
yeSPxaJ1vM/9VFaZVidqaJHrzdTIZ/2vBR4nUeT7tU2u0jupsFZIkgqYnDpbbPU8INzHEWsObG42
FA2qG2MWrtxYjUD8qwkZAooxVmWHwYLGO2RGwH6gJZJZSLcC9N5DtQ09OE0FRWyBeFbNEmnizHEF
bMO3kLSaWprCSIVVpbVzUSUKJd9ABgL7MYZSeUmm4lwpcAAODnNu8+zM9TjBNaSEn4M2Nf3drxX4
px+3f8H9w4XFJvy5hp1H/jskqbYMs8z10vmv5W7gb2DLNXRrneLbbntZYHOZTZUT8wLKK2JeCO/T
GIWD7iU7uJ1vclV6J25Rl+5Cs3YbdgP/aLE7l9/hWiyXs6qKlOKpKy1TkcbA0M6a7m3eTM/TRFav
YKVqKqc6rr9hCNYlC6D56vA6gaydDD2Ap8yprhIrrYlevRT/swxtzvqjuXy9wa89+tvmimecdmd2
aPS79VvL4ZYV60fPeRmoVjgdhDlgC5LI3IQqWXXkrqiiuyKXYxGoB1LGymV4QhUpxwCUv31D/pAU
ltqGn0FahsPcb8ZNBrKRuT1Jv0CzOW5H99sMiVoehNjevGhrBMDvu+83B2I2g0ZiMkThmA6Kbv9w
Nx/2EeqcqRm8scWf/xaaqmfSMoZ368RUIQEpS8FSP3X8/z9BrSSW7q7OfZyhw/eOan/OWgh36+zS
FsiPSkdL/4gd9IipN4JxgE1mhtpw9ip7mDvXN9cSIh0DSxT0nEOfEQETweIqF9v2GlDGW0lmQ2VF
ggQXj+1J3UgaAx3iSNAgZVqxjxWIEW4oLM2vTvVZtLALeYb9h62u7r82Q6YsbPRdkrls+4Rv21xW
Hq8C84YgGMC1rYKdSOW/gbQ0k/TsbbaQPy9QCHW7/g4LtBEFwvARmrjuvcsuX7xmITZQ+P1BMC+K
DL0YvIH4BUioYT+OgURRRv6XzEw2TZ+VPSLRiketx+LPhX3BecdJQQ+rECUmiYcEcGpTyFJocnBl
VMmMjRM9MO6zIVB/WTq3+bfc5rqfL8aacszK3uh7FEAygFSNjcVm6zRMxgDlG+I60yD0BK4GLHlV
idwnKZbp3L/iqn3E4RHwDXT6JiEO68Of4VhN9oOgz2WhXwaA5Nbm5ZdszXgtkrzbz9vCP/75nzQv
CeGZza25ckwn3EOQgJYPo2ikW4Gf9uJKp+DaXis5hsKqMgKqHeS+B7LlomfNn7jA3TOoMYDagB4v
Zh1tNmMyypdyGEdfRGAxiWg0VugCs50jr3DshJOuea3ZKn6IvfvX2ghTUqjgsrd10cLWXHQEagNg
Gel22A5Vc1ebWteH6hUR3/lDWz9lJB0S3pgP/QCr/bc4dXKhnhEcDhHkBM4fAau1SwMJGe7kavxf
kN7tu0mInwWCo6K3Z25YaeAL3RiZ4D3w6kO2AiMC3mHDLDejpUOJFNRCSEH9+PTCjNHvotsqgsSO
KtO5L99SJ7/gh4rjyTOpGMgry+XCNQ+Hr6oTi/bH4bLTSI3Me6g4lfdv39vlsGUwHDC2ioqPU40s
n7ZydyGbHKr9z+rtAJM0szEoZR6MHuWlhqzCG6ead6Gspg1ZEHKhYsMgNwoje3J3rjx4kSgDEIqy
TlpkgT1wRU3J1pG0a3mpX80LPqvCG0kt9rT1zPum8uTPnY3dlP8nM91YCCoBOIy8fL4/8CTzjlN0
SJ0d01lXv1P2EwHeVZ22ltlRya+NE43S+EI5zM5XQjSo3mKdBJLggT6cLDrf5C9+FGg5Dz+3gjoh
uA/pJjtsvjSvFGq++dwvRnJLy4KjTK/FEc1QUrCU6Ly/oEoxAXANfZg2KoooZN4iI+bJiyPKy6QU
OtYwTt4mmjr29SJ2uYuvjhvjvhlSAPfRfdk4hH65e5tZIQMWJFtJ3+RXzc8shHGBrJOyS6C/qNUA
bd9H/utzpY32NDAARyRqsUMuJVdvvigLVNv8clOV06KyzVOdf7uzqar0O6Gde2UsLo8+WRNXf7MM
+TcDGXlgWNZNyv7kOvFhsWdh/Dd5mJAcRUvKO064dA9XS72fTiukUCFkV4JniunuxqzPcIg0KwxH
0CEIO7sW+mwy99+tm1S2HaxETnrshXtMAQqndryxIZFwtB/ErROwGj4z4ucXWIoQVe35llwH7Z5Q
FblEJiab8Ry7wFWstJU1XC1zDgQVEXiBLSpdTFIz9r9yvWkR+m9Ay6rUKWgoPUZbDI7M0MLhhbAc
VcEthPwPqg5knfZxFkFruWbBGnRe7wR5hFVr/q618+Px/BT7Et1u0ysTuy/Arvg+RBbIgQmSniEv
62nm6NooObYtE9bSfxXw5SRKrY2hW/iMW32UuUXC8bu7gjT7c6+YZi7qgea5diuwCMo3+dZDEXSO
745F8ICYb/QOyr654NITdph7IUxxcy6ZbB/TEoD74Vus0tdm1EitZtmQH7zojnWuW+SuLUCKlJ6q
YExRVGFu9TPlF1oUx/AFK0I7vAJVysfCQjK+mCduL4TWaA8emDwY132bqfCoPEwnE4bl8t8QiQ7+
bpiT/iLONDVb2VEtHmT9cErNbxsCiTwVhV/50kcSgtqLKUF/hMXWFZHFVrVS8bmRPeLa+yczRy/P
NReY43c2vHbtqljlQry1JimYzikqjJUycUrzboQCDue/nDCNm2aLS1X1bQ8cZqmPJqXDUINqoEjp
6goa0fNp680AUyz0D2K5hUZ9AfA/ZQjMgkjReWqjtHF1Iwfz9p7Yd1Gy0zBOp0vu3qy0Q5Kxm+RR
zcQg8LC3x2QLhxZAjnBy/oDfw8jkihemB06ZBfifkhp8VQd7B/BGtiMf2ocfV7PxfD0a7WQqXLus
z3xH2sofSFKy1ezEYoxrHCjO+JIq44lEK3ddC83z/Upr/tmCiftM1210Xtf9SF+icAWzgoPlNHpS
8rCZa9Q4uSNCwxL5ScpmIvzXn4NBVQjIJRTVWfqxRfqTYGybbiSXVFEkRBW8MeuD810AanWO+6hH
YPqDTryXFyIqqJ2JjkF8rFuNQt802WcuA2P5aIoBsrgi62um/tRXW1XkDk+1b9GfRnVQTKw2bqFl
nVhvooLxp6onMLS5S0sHm8WE5DcHxWCxQ6sIjcJfS2vnhF+t82kk4YIS+xbTXIclwi7qlPqaVD7Z
20BeLQd5irEg/qe01Det7yWmkmwbG+L46IJSFUZlS49VONI0l9PdjcB5qWw4KNaNHILFVAZWoSeU
M6aUVn+CFzPCoW+oB5FSbWfSBU+Z17Lal63ADU34R2cUmT59m8/bFZQ+B8UEpXTCx+r6hOKJApDl
6dSWwbOWiODBFFGAfUvduspEByHQtm9hJTCy1gWEEf3NIqvQnile/SUpwVAnphuGx+CQeKMRdd/e
fhKELL4UQaVrF7+sQW/QgaqzOH/8a69GlDtU4O0otya736MLh9JcRoQs0x59ogHL8hVjZzaw12tb
Bnz6jcDwZ5adLw/HjEfDR3qDF9gdFIlcDh7FR78nTFs39uJG2oAlXx+woYYTwpKvAR0j5jTRkZWv
rExCKZ1+MUPo9zYPtN8Ks+JRz00vF0wFRz3INtbKZ59sJVf2RbHAo4bVk7sy6Fc3qHf3jqZAgby6
9EVLBgFghHMuI0lRpyzQ+7OISKcWcRwuq4tSBCeFLQqB0joqI0zUeuozj12AqKnSR8dtUewVIEej
VpQjg+5bQywFOWYxKluLPWHsCw59UqTigtfFLdfBKhN2JldBeBUPdhdfau3ZphE/eCcoFvSdFT6a
hcgifFg/SUiSLt42+osTDZvfnQh0iLIHT0X39MB1W0XHKhXy5b59d4PyK5hWwqAJjoCRO8URYNZq
2ZGhyI5QpTqIxyv9xWnC0kZYe/fTih5nNnil1fYa2LefWZ6jZ5LEJp2pMcy1YHd4A4tTA0J/Vrg+
jJX5h+QPxbiaJZ01uW8W7hJbREA7p6gUbmC2pmNsAl5DuNx3OEceAYqsM4kU6UKjVotS62XUxsMD
pdpQhZGVL0UOPjJFMW5JOCT5btd8az7KSlrCIuLvLxKuDviYgDTQdkg96nLz/Sd7h4Axxtj6ZGrv
ao0VAk78n3TEAq7HUP1isFZJnpItUhO5UOV8nHKuz6Yn1bSsgzMSFJpi3HywdmY055f+FrmJn3NB
Wl5hvjqDErZa6J0pGb5HK8u7gzlyU/hUCgFzWZh7oJvo2FzTSIFM3YKGVn0rRfc0ByYpTnWLg2/E
VL7BzYgFm+tvx0WJSw/TT7tVywqcyJoMp0QeNKqTW6aqdUd/OCrM20McHFxdpYrrTMZhWXIlXlYV
smw8Wp6em01zQtw7+yshEieYiKKaLAxiOFDOnWZ+FmkJS4ICJ54EeYlRCDpASQR3ZjZ6nB3bPWyH
aeu01e7jm7Aie1hVwYmbELMskGRR8MqSUMa+vQncPCIllKkuFmgSkT2d29Fh1O5ubkk3HmIhaTvn
Sj9IYdQOvVbMItGJV7sLdh7h1mOwMlavlTe/CQpBLrCNxDJGX8K/XPKz393Iy9pN8Na00SSgYL3G
Qbw6+hWsOMEINgsorcDXSeWAPESkTqtK8GYEuKzkQlvmi9GRj2Lubs6m2nnWIyK44AfZ/JQppdij
E2ZOBoMx7zMbrRbuJ8lDVKSpAB1B/y6j9WeEvphCGKuoIAXM/8WoqifopKhujq39Mk1M9U/UM7X4
Qp1hgfVXl1cRQQkKMKLmC9L+qRmTEFGN9mA2QafCb6bPA9C1w5BeEQGDvKbXdN6VRkG0lHChnMcA
BlK42OMGklRqexncu8IS99r+sknqpDa++p+4wNBJnUmuwsYiQ3ZmfVpAQ1oMsN3XHdhnb28wPQ+A
jLDAPyiw3euIYr23S14GPcnYrFuQJC6qOHFRJby3U1xJv3jJk3uNv8f0ujqWe5qPjkTy8eag2h/A
GrHLppHw8GLxHJ3h//caR2SiTnE/0sEF9ZglYHV7gLO050uZbBwBSp/qyuoe92ykHfgGW51SZS6h
5dY47cHT+avvr+mD//qOs1KN//osZlal/kiGQgkquTYeOTuReZoNvLDFbtrFD51rR469+eHWJVTt
zjbzlA7Erk9auO3X0dCzp1oSF+2lX7gjduEOJk1zTW9Uh1XwW1dIXWGBCWzilmpMJblY/feXjnEC
xiJIZOaTJNkAQGiUSKLanfW0HwlvYnTHDyntzsQEfYAbHFhgegXOvWE6+FibdYshOPoz+Xtp563M
yn8Qn+9BOH7P/LqMG8iADX0TqC2j/11tPJX1JRbTNuN6jD5msoNzkSu+miSQ6hqhTVgQAiYeHB+s
sTN4lCJc9z5CViZfSZKvqwf1T/RIv1rNjhJy7Tn0+JSdQuXeDJ+Ai/l3D+SZHWdh9TFr2V7M2r17
y3T92VqROcml3wkbHHSkROeBi/r0OkRKkyOqOzqJVhiXto+qjVpFftEQBWna5j7OxrKwt1GLCYbf
WfC9lpgrexySAq6bo7WnRapriglNhMOAxV7lCvZpOno/8ED0RjbsHFy2JbkWDKki0uJMCR6omhbO
PdlDzUeYyguERcimqh6ciacHy2iI5dTF4dqmeltlGgsXd8yUzTNSHnB+C0NoTxah9DsYXqVdfuAf
9UopkcQzbjrKTqjdg7DBWdUPYVn0YFej390jqfAivg1xEZdrlctdt7nYQcv5EPXBiFb8XD6IoTYl
n3Ol9iZDdz5nPY3fjPTs8w9KIrwp+o10hcOtRK325UnaPHbXgLNv9wAGQQaRloz1/AE4hvI5EEmX
2bMsw2oYXvPHEMzzZcpjDQ1mbl6KFl7bLuvHMM0Y57UWc08hA1HHtlcl7yeGqKeg66kULPRLG8rn
nV6bBPmydqVbST0G5dTOoiDVq71kCn3k1ba2OLniRSxhc2SJpSr+5MvyUhBY92ax3J3CZnWWYQ/i
Ca8gJnECsXWEQ2pqoE3Na0ZvnhrB+DXooHOheGi3od5KAelwZRLukPoj/c+5yjHkIC8F9E7RkjvX
90AZl3FIbsJ6RcGwO4trE6hbmm3tdK7lKs5lk7RUT7AxOKvopJAABlN0CSbA7H7iZaOMUyqiT3HS
W0GB2C0/RE/YwbaV/zWTO5EO3JFnsQEFndL8pUqaHO0ZSUYGtcoHl/6q4146G/nm6OpzupwaZdUF
bEZRkmghuC9TV+OxK6BddfGcMaFSO2SvHKHns2Vc0sMr6BLtLVqm12LxjBjGdkgjXq8b2Ir6nSIR
kEF9staN+43e89PqOY/3F9TQILQzfxupqI1TsTQpHOW3zlajCv34hGmW58qqHdPuFDacq+yCNLq7
zAu5z98m4SS4nEc9V3ixZMfHI96qgQRnpsdgbUZFt4rSyVnEYgylod96RqbX2SfB/kPVgfSNqi4C
dc9t7+aR/ZnsK17G9NpU1kJKX9Lw+d1NIuN7dx5N5sLmDN+7fDkqDVNkrjqyg32S+RESKsk7hltc
Hrmrqb08Yi9o4VbdpWYrufydYomB0i4b4MjdH81msbh/SjDUs4cxoDeIQAJ4bUjtPgPpd5whB3lz
zmhRAcN0pYz/9qV8eMiRZ68YiWL4oOoq+mnpz66oL3xZBlDxwogZZIoFNtpaI/yNexxMP6DR57qn
3ridXbY3LSKfB+f3uNtVEgWVwcy3zznDK+dHnIzQBaDWQS3aIfFlbK8MxXy2ry33Tbv/qEZsKJrg
NWxlTcfNpm9UPlHId9EC72AnEYqKP1v+7KfsHnBcm2evZANhOyh+kIf86HBkNpjsaiv5bsH1mu0A
RRKKtpCXBKuMOeiG69nT36mQnnZj+vEyur0zAwRWYFSbyguvVAv4HmjC2Gho4oOSI3WWG5o10klb
+Yt9/8UbNv67Zcq7R4V4rAKmLXx9DdUh6d/YhNRuy0bwXN/Vu2y9DY2HortPInKUgSQGYrwRX6DY
qZ8P1XK8qr5bpoCmysIMaw0Rn7XzkO3lIxJtEREbjolb6GZJDFcuFFalDtp+Pa7ZDIdJNmQ69MZc
X1PZMTpjuaj6Hi98melQHS2wb5Cl0mouos4G+XJT6oKJxnKuiT3jpDoYw0AM8ZwlIwOvQ2o+l4nB
fFYOg2qlxhDm9zSKqO1FfPdE3qFVWrJL5h/1CPaXvKP2rfmrKdXpiq5xI/Ijou0EWUw9wpTjvpgJ
emYxwHv1kjKtG0aO2r9IQDi0uI/Ufs22EApmGC4FCf8h8Iis+UmpR1HUbDHve8QA71LMny6g2T03
NcLgsiAyCjF9t7ZZsegQbvwD2oZl0Gi1DB7YQPefbuRkoVj4TKsWAOiIYg4JRgCm7rrC6MZl/VU/
bhjdnIGWwFv/fguBaYeaiOvhiKGbLfrVNuTyFeCatYDqcsGGJ3TkqS+VYJM04uukIEYZ70JSUknN
ihfCFaG9FiBnV/GnhqyGKVsJLmTrOVhAkVzGjoYcsnQO1tB6E1yU265NX9RFzjqwROuxTKVg7ATP
WzvL3RZiRDTUW53/QMQXw1wRQ/yLamEBFQHnrpCXyyHU5F1BOmJXvINRJgpDDLJNIVMp0MHIZMTs
/UAOu6JqzJIhV/ABrOzp8YgFX9XFRyb0OJ3weN6vhtDmObYYHFVw5gs/kolVIitOOirByRBkU5x3
DOKppXbWVfM3Top8Bu0KTcNracB7EgJ2yxjsk4TMqxKce7pnYe9oCZciGtCMaF6Sib/AgDpEf0n9
ODN+0JJHs4jxDKcy+HE2LlOtCNO10oiLlfnPfiCbMcG0Rb76Lot7qhP5czMU5pITBc6fGSVQIFnv
/6HXtLpp7RpaJ8ejHW4HOSYuU47U7bYxX3/u5DB4Um8H2n6WbKzqwpkICSExQZ3h7XKg7st9wlC0
4XtyZnlzSyQTzkiJdasE7k1yHsB5Ehyi9d3uo4ShEI/34aHLg1+znZz/I3NO0QukQm3hM8Q8tUM2
TVWSoL5fJxOTjMkyv8GXso0IuqCUugA5ccpxVNW3LqXYrj1unt8KYTeGFJNQCxvlV6e6eoprlNHI
THm4ECA1ag/Wp7YR5RiJQDNQigonC5+K+GFTdRSTKEev/L9jICJu0HLeoTJu0mB3IjVvbZb7OqSh
6x6tBOrIa9t6I86iz/72iA6ujcD9esfOMtEsex1GcIuBjBgLvWkdJHqxFSoKYpT3zZ9PZPuvv7+y
Lp8qabRQMGtmMUAxCIwj8dYS6buXAD7eEHjlLEmtF9g9WYJ5hNFcTr+GOT2enllUP5CZFwtqgg3B
8ui3LLUOtzdgu0+utRUP1+5itXLemgAP/MmQtkRo9tqZNFcVeIdTLoaxhfZIKWNl3ZkIq+9XS9ai
elGUIZX4GTDcLFuXUkrzaH993ZUih66bNvq0spf9yAy33pKdrelmdUyO8noqmHyHBv2EuSkcMYUC
qC9vMe5OVjpl7WN7FDsPc8i3stYlsVgN+x/UucuheppfZBxg4Ma3pxCEM78ewX7Lvr0yt6yg25CW
BRC0b06/jVMVB87eynAIlcVnT74YG4An8Lnpoj2+ZiYo8vSZ6PV2C0zzKeRlN6yuVDnwS0xv2FB1
YNfAUDyXYijuPfSgxID3LXzXTzpuiHI5GvRNVUY5iww1zsGmvCi6GNPRgs7F//3+bOqOYuHxnrvM
zWi51TMjMZoXP8mBKWOdgr3Kmb5eg4om1gWvSm7REWEpSVA8HkksWTe0N9XfkVSCTbmgjROAYGAE
Fsmgromqer+OicYiWIT8IDPVWCFYn6AhfBh/XmCLTMFByTchGrTvuckut+L8xVD9NoZxr+sCmSMF
Z+58IqMPskSuoJv+KSxo+s3uX0SrLo9/+vWd1dWptUprafPsxWcfCiU9O4fn50hyEZYme4/cQpfG
RTQSQyusMol1bVqNSGDLFnZsE+ai3z7q0/s3+1pfAPvchGTrYZJjuTwKXI9+IwdSO7S+ZRuBL1zv
J2vfz2pL0+dWbQ77GATHhmCl1iGGsGShUSWsrMV72vA6um4z1/pmmM3Mld+dc+6ERi6IrJ3u8p+5
cUvazSy66YVvgyI6r5owtJ4pvwYVyGmapDakFUBadMEEq6JBJg83CXX3krQWEiL/bYaKDf92fK03
Q98Til9X3SDg/q+TqJ9M8X71SurkbRYpILnLLmlxc64t0FFdhTwpQVZSNU429IUIH60jGgMTGOxd
HWq0fPCKgmjNerM+Txq1FWRJxBWGgw2crAkzYboMo607ZSCipWnkr9qfOqdlMJx1MD8V12KJF05r
JPVsRh64+LhsFfHv4DTSLWygHl19RvXyZCKAL/QE9lH/EBkLVbSS/t2IRvJEWJlxIlWoXEd7I70u
loj0qKSuc5Y0Vb4IzXMveM4GF49Dz804aspKCJ2UqGNwCEUByw16Vfuvgb3s/9Nig47ntdUAn2Zk
d1yZ+ENyWRnYtEWXsI8b7zQkr+8WRRSyYULFKsHssd9huWQngkiyTkvcRHi/l5ICfneZqbUspNTa
u+uDTsWJ0eFJsjivfSTghVObqsTfE6KSX9oCAeOD3Mei5CaSJB84l+FD9KqwxjhgmTvLa5vNrL4D
QB+CWztMs8/Xq9ejUrO7EVaM3wyfiv/xW+zEPC/bAGEPV6Mr3lPTvsypw1/Nc29aHfDM8umnsJTd
pmJ0MsTPIP1mKHo9plP3mLHVIA/5F/h+cLvs4kgNio6wdShZ8UnSAhnfWwnPy8f2uludnzAJobYd
8cQUBmbNm0GyslGfYf79Z9ZXI4lm/WGgKxBv6nJWrquJAZnV3rUH+N5ewu9Gf7TsRJzuM+aFKle/
JDtozDvrfXoH49VSMoeyKWcc1Tu04VoRJaaTgmGiS+rMdJ45sqv4WcMJcVCLKN6HFTaaVzb4c84n
bB588OQbpbXzCVoQhcQ+XCtd3RfY9hGs1ai54DfQoiX+2/AfSRX2yrnVQq63nI6VdYrWEe/yJLXx
+zpw+BDVj+0gqCWD6ymQHFItZh+9Fs2t9ABNib2grIbeaAKhinEKn0kFLbNIG/FVejr3G0s6W7WK
LEfCm1er4TVRN22qsCXUMu8yYmdIMxFrSUIdrdKa5h5D4Se3ZQ/P1W76wIfhZsAwzuU01JZVHmhj
wLb3WrnbEneVjvO4H/EaUsy6M9errgEl1JDM2DMJqyqBJxrTp7EKoiVq7TPyQm/VbHjDpolLO14Y
JEKv+iK/vjkLVz0O7PwLjrNU/J+9/BNp376n/t5mcW6TsCyE8ySCPubOjhQ6X3FMLCfqWZaiLhX9
vzTUWYNcPPNdWjOZLSOuHAkTfpneNBg0Yo4Lt4K4k0aL8GsqlTWetTHpEcZJB+UymatMHeIVfFav
pJG6SqVZ8+JYVoCQ9GusaNfIZqvNFL1L0gaUI4hq6BuM1VnFil9v2kqv8+y7K0ycKwsG5ikikolz
nYPtLNmcwo7mS8i7krSX+69FP4EFnE69umVYBqaw9Fc+JW2ue+5pBCWgkS/t3J7aMaywXE6WbaGD
PhbhwuwmIHrg4mW4bajadj+hPnFGioEA2iwsOLHb+dTLeFMhAhfz4u3Hl0DlvHLVZYZgRVgvbzGz
iZwHHuk/CGjLe1NUjPwntlAd85QOIaPhi8Yj/qMaQvYMDgZR/sg6ES0OTA2U2l0sHXCBJBp3Ju/b
fNzsDKYNC6DMtDJbUxtOdr+0p+i2m8muKhH+8jFEaqU7/QPKLyYSp5mcEue3FodHRZVL0civjony
JtDGfpIeRlK74q3QU2uiuOEQO8pbk92UOlsOk1WlXh25l3Gsl4U7GdRlZewMbocmXDGe30dggdX0
omDrKVp0k5XfQaxggQkyP6CU8TeozyrR1ZeUivcaaiuf5OnlbbHXQtFwtNIGzZj8BXAqB1v64Wdw
EhZwvw/VJF/ZBdfTNtwnL/lxmhs6YLigihx6hM2guTnWIe6UrNPCpBtJuUu/NFLmxfSZlEBC0vf+
SOM+iZqsmOTA1BoExAXMjTTFx7u7nR/IaJVjdGyZAqsp4re/xSZ6Iz0lHPgB2VEqJLK9k5jVK3r4
CxQJzfps7rDqNeuDkfax+FFjdeUkbC+Znf3xgZEM7ytJDZbLXCr81g3WtJnFT5lBv3aUUfPbBhTs
a1/TB617fRIWDYUcftOIkRH5IG1WRxZxG7cG25BevJdFLgTvzzjWR+qojgWbecIMY+GbWr/5ZfFF
bM+gl6yZ44h4nrINZUcZ7Y6knf/u6aV9Mlv1stoIarTNMDxg/Iav66R9LHIQ9kuVdAy/qEN9x+Qv
SZyHoBNN3CAcfinbPVbSuNG/n8PzQVIkzdt66bmUjYEplPqbdEHCXlw9Kakaifmy8Hm8XRmecj4e
iVkAasefXACEFpPgoGeWHvZ6ecYL6ILHZLtctE4S+Y4Ygt+BgrXHEaCgtz6OrWnKJ8YCvIm7uwD4
0Z/0e+IGZ9iBHtXg7qMvGYUELXv+Jn2WA/JXioitLAiZGoHw+wWd6oLlwUjzZ0W1ehnAR1RM5ymE
IcuBHaJTfDYGmtrDiQ8xvQFAu3VSOZ+nJtF2xlei2xtVn8HOc+kRKXSqhmiv20eYM5anmvfo6jbY
7VmJ4di7KYGvjWunenuBk/oU4VWlNAMcyLj6GaWVbHnBKan7INzhKtPooYkn9mahCmv3o1a911AQ
WN0C3ZR4q4y41s1CLBChNjcGVSgG4w1SrsxQWss+x+dVYPW6jvdVYaPqIWqEVuqK7d8wbubBo+xA
EYYSWnbVNucWgUo7EA8Rgk4QFvI+LtsIxDDev4JCHcCOqlonQh36L5EO8oeoDnFIG+pedU2dc6Ty
bFgLILggL28ztvIJNqnioLpPne26LROW30MT6NF+b3Q2/SBA8OjwCU0sa9jwi4lvWB0TMgmv+sDX
v0qOBJisxgKxbQulFvcr3HNbNVMl3iBAxd1RgjByBotvmyKXY3ufc2Jh6pkVt+ozLVFxswJDSgMf
+sUPlZKyuPd3h1l2yQg03NE72DFrVQ2unAldmWK0IQJ7IeNE6+q2IyhLHFtufm89BSUyDC65hLLj
6LWmzUk1wMMFzn0Off6grD3JmSGLrzHCn/nIsUaRi+TdXYc8dZjYf0oCssIKvmtgbS+uu9IoB2Yl
2kfeDVBIgf97RPJFrAeP+wS+7jNo+N2W1eBolsgrm4TSNmoV4/W/akTHFURoOfUPOmuHDnPJmcas
cymQECcrkk0rdUweRcnPRQdwp25zqCl90Xm8wy9L3bK8+FLoHXpHS9m65iq0HD2MvyBz4M7uaGM8
hxT47h/60FFTc5EDyfsQh+aNw7NnHtmyLL6hsDNFwSfI/4LjpaOBfcAGjPFkBomlr9cHKhd+NaWZ
dYEQOa16fDV4zH+u/MpsRffSccqU5Vgdj/4luGaCwL6QQDuoxicuxGIrWyX2kW30FKnRX9T93XfK
o1StKm0qOU5FsOI4HVxk3NAxjwYJy+ikVuOwOct3Z1MG7jm5GkAXC/WVOsKocVE8tVaGp4fKLmvP
+wgGr+MYVzVrsPAsZvFIWb0dHsMMm/N3swKsXnf7ZVlpKKyGp3QpeHu3Is1lri/c3TP85pYHJEaf
88I3FH750d6lMepTWYrIIXmFDozAl9o9UV7Pn4z5pf+IV+uqkozWDUrC7BYJBrpcBgKkH2QnEQDa
Ch2M1U8UABtMitcXP8kVY16PLbl/6T5nzFw4WAVKRvv2XPdaVAhBLa92o7OqlL8GiNyWT8jPWMAw
7Mz18qbY2a7ZSmULf7nqOIm4MpnBjCsV5ubKFI/gE3hzOoZOsKTtVwQeIwrOxSSKiFRM3ToRkfeO
Oif9iz+jKqqGLcuge+lyyHvZA0HgC1VFfu+0xU7P2cVIJWjJaq18b+koPlSVFB+1HRLcsttmuQqj
Sbv7AYQNaOTCb7UW2pEgT/jPsb8KM3k+NByDKE7L/UbLL265u4h4jmtyX9tCtVTE0Xy6dPOMaTZw
lmwvGjxCk3gvgPDHHZsZFM67wrQAuwVJIGaq1foaOBR8b2rmcCR+iJtDqsV2MSdfFm+CIVnxHoBo
84IDDNMi3BFv2fFEgDadSZ1Jo1b2Y3rzqktR0P/OXe6qWbhRCWBXkmDcExGaPRTrQkD8YL02u6SP
o5s/L8vU0XhjQW4s3Z/EjIp337NNIWBE0mL2WrTbwePAaHKca0dzpwF/bCFubIacEcyl2sxuhD0o
GLeuBV5O7MYLFi2oVDz0877IFBs8Qzw7zvqnqeY9elfU7mRaoZXfQnJO5mM8AWLuWi/JgWSo/zS7
C1UxZbSgG7UiE+R2P5KAJTN+d6XSvqcutLEIOSSqKEUACSEFuld7yRYQAcK6ptEEouxmMuxLfX93
KWB5EZhyKi6ckmlXll6pD5Q7p0qI4a3xUuB22oIEwFuCwIp8uJpchMO8bWYplJTAjenQdq/aluA6
s2kd7a3RGhzAJbmUBQrmHXf0NmpNs51Yga25jm2LxAw6vqxDyFx5m0qc+I8ycAxpW8ll1YyLpctk
D3PbUXmwJohxY1PtpdlngF8Ge8tnjKVfzICcQ4DvMIr7xN+0sJy02Uji8j4dpZUWUhDpifCIvj7/
3uiya7MO6EnIiR9DZZBsZchSn9xFDSooFfO9JCQPxJK+YoFacx74R0yh0gpPWw6Bor9Sk5hf1TK1
J5NFFm3RnIr53FwbwtziwNRnzw0re4eoN7i7Tqe8GLlMeXiCzNkOnocJQ8oGY/kxh2yCrtNK9cNV
Qm1T46zKQmai2dh0HdaJr3lAhcCpdL7gMjakk7/c+4ve1yGCSc62JnF00BDK+v4K7vA7KJp4+YzS
14j+tzXbjaMlGgcrBMm0AqSt8F7WxCFARZn3Nk9Ib5Tngaa0RLd3y8fSyPkBmSxYvR9A55RHfb9O
HpmgJJo259SCuJ8bKP9IkDSIHoGKlOnLOaIyq1kzEbnMg7Tqz3zMcdzTVak5o+qKO5r+ZehVyqzs
sEuO8XE1uaLzw4sBhehD5I8D4v+wEIplcBb7wOtv0GX9AmEDmzGZPGVCiS6Vyyl/oXthbGqJOx+c
JtE7vOpW+eN+G0pDF3Tyk8aGVbVX3EecMlxlqiEEvZRiqbl9NRwKjIKcwGuJ0mGkCqvFFc3bLWr8
RsX34iHxAcXjmuJINXUaWXJpche9lTIm9K0YtNwSJiZOziYHh2FcQKwa1k6Q+2o7eJHkFUMDzPJj
lTt4tQ4kAY/Mx1VkJI74Ne42sZwtgOXNh9rEwUQ8QWaNUZFJzTjgLw8kF575N+7DzYSZq8LFFV75
tVvxCVVyrpDQZF/cYixxNogxWcFp7/gZtg+oArOfCG6jdlAxljtfO973INNl7/j29pfDXcaf0N1P
JtabTROIFba6xU9CGR6vqdafXBG+LRHjQep967Xnyh4IRBhEfoRI1v1wtQPphFzwmMcctFYkzzQo
mo1hX34MMidu+qHhwVSiXpRnSJClaFEyS4nWpyhr4dqqrm7zQrPtIGElsgVQSfmiUo6jzjwdR6r4
/7CsQjfYxQWG7DlXUIXoe6AZyUt4HBo6My8htOgMof+imoy3HnM3C9f4oGR6agMqXp94hbngxomK
abnLuoVwsjCJIcm6jaQ+PbxO1GEwBe2AHXYA/MRKBaI5k+Fo2Hrk7Lp9yXrSZIF31oMGIAjWWDVK
YIOL8l/CHbwASscPsGeXxES6vtry30XGiqFq6jWihrwTBHJJXCJYBxEKDBAv15BbgQ4vHQYy31pS
Tovq+STilwDnSCJU4t3R1hEKgf8k+VLTa0SHEScOUNuTVO2DBaLHm9Uj35G6KIXPPOLugjbcCyF/
9hmH9i8HqwN8v9nfhKZLnfHhxL5Fg5QXsTVXnioWrc1j61UO9PIcbeAJit5wvqdQoeVsAJGJfdc5
jCvtISU3uJ+eaUo9Fq54IorUy/atOOagdAcbJqeqj2VaiX3ukKnZySXjhmP2gxtrz9eHQK+ZD1RX
82LlOknu2ep5pCZ8PwM9bnpL7M8mDRwumP8y+zffAIedDF0XP6M4454weLrMoVZ2VpBo7JCuaDe2
p6mmhPd9k26IZWytdkmw01OwDrPFRkbSuS5gFLq659lub6Ef17Ivu5tqqqm1i3fHh2JOmpfq16Ax
5DP7L5Sxg43jHH3FL1VJYt13Tx+8l/5bTJ92Bh+WgsINxI3EY+T2dk0uxBvOihUxSIjxgwdCJSZz
HvyBDEMR7sUutU8clxdYTBJq8oNieROyQlLWiuqXFMOqbdKqntCZWJ500sdgsTIdtB6/G48AD2qQ
j5QsgWcYxhORIyg1c3qymN3WZCtZegyjFHhaZJoaMWOM17Ry0FYYbAmXGxToiQvaLw3BC/JEQplZ
6Q7uz5twA+mZzbicCr4YVRPSDvn9ZpFTnsKiJsURI7iCRvJb2kKIKBexerdz7vYJAISovS63+Lc2
RGZweFxpVmcl0WEPY3C8ksloZoMTSnCNpJB1PU5v4g4hL3x1d5DGN5Jcd9hh0+emhQCKN5IdfBCq
aYX3SFeymjkakeSzg3bP5w9msS8J19dgkmWdDD7f/uf/kVf2geDxKCHLMfYWBHPp04lb75/1aYme
+hQ39H8UkmOOVeq7/74iaHsAD8hV7XmEgGG/oux0EsGqI4w+ZJQ+mjQ1fqYrT5IOhBr+meJ8zBOB
oSCjwNB23anwwIXSrxv63tETd6O5PKsL3WljyBJRXquTpGKjalFRqIUoCWmSYcV5RjtFrcoBK1Ay
5mPcP2/W59tcUQN/WgHIgs86UDOyuHg0TcYxQ3K+S14JsKN8yfD8TPi1rGL+BmZc2JUAAtvd7N3j
+4uDmV5NDYNZ2r5gNY1LWVRb2r04Fgp9EnY7QTD/2HGO05vLavcVdho+z/E4ti9t21y8y82+XvDj
n709Uo492xzxqmkycE0suQSD+yZpxVML3gZhHFva4oupSKx/RTg4Mn13JqBo1whxDCb1DxxpJXLQ
Sfy6n78yRFu0ink7W50p8yxNHbBFlifpb2+jGxQthGWhhOv6Bv3bTkuEAcNQyslZSUK4dIHFu+bi
7aOSomj8mQLccY8nWDzqruYDIfVtto5TKUobhmS8cK8+lsUlS3c09yIUkF5tLGZcYAIOGPimwXsd
8WC3VNKJOvx8FK7G1nKSpy4SrBMyGTH1MzaQFislKTJEBopJEzW2LK9jnG6X1XKP9R0MzdVI8VTo
8PdXSNASzyEXh4Q3EyeCVy0h+WE+hyEap5BPLQ1rUIsM97YjJkcv54a0mBHRpeSJ4B1JsaXlu83w
zX0STtNxUMAQe8u/M91XWcqJHdf3HFt5MI9xbF0ahTZcwYTKEgAAaRlfCkKWVdxjrtpaH5aDJErT
14X4h6VOcirAMhA/lYBD2Iu9dq6mOoAXTeyBCmRgLlCRMG744RQJF8+DDyJTvDSEERGWI8yNWvZC
QjxMhfE+LdvPei3th9+oHrzaMXB8rjCyYOqAXPK6iTTgl9ODXmeEJotQQea+lPZ7QnNO5vukniQQ
vNgb+awBa/9ccJMh4aVunI6G37kM22AhJIGbY6THvKtnMlt9X8gDBjGN6t12BXDztCx9N67q6TaI
1BStZ4emlAWzJZaG+058TgEugo8m+vGqZ6KAkyu+F6ufgPQRTzju6//Nowtgb6qF9nA5MSp36nPA
my1OIxO//7AtG1s929YLoWmommhqim4wEj6Xr0DRPeSOG3qtBJHO0LtYOqe+DCMjZQj62XgRcPz6
dQjsN5Qz+j2M6vDY+sQZtYMDHhVUFft48iGGhptIZVlOg5CRC6okk4dYREov3G/91LU8uhVYGEjW
70DC8CVqxWGcgxr5q2JKfYkSFjZy+l6JMUZattRN/XalRAUz2eaFB9Y+d3AWap4TU0mtZC61mDzw
9CRIvzUgwQLFrF5JrX3FHYPFdY8MiU352qN9+VLPYvqqvAV6ZNfL501HDXqYDibHar2l3gxVTvWt
5CRhZP5u9/idiJaR7e8ud9t941pT7QS0nExFJXafN0eneWE3SKXDpbOAKerv43zRXDJay9SFp1Tp
4/d1fcPJZEDzGlaltV3k+JjN0jnxvwvCgaQ+d0mbhYJC2hoRavj7G9iozwEH1dIYO+S1w83LrnaQ
j19R4q7lP9kIVpDcF+m6c59Cp0qhpH9eeGNX/zGhudfOdellDCGDo6F3I3g1XU1Z1guxI7e3I6R6
5jOTY6EZCwgknrtpYHUXRmwl9Mnq47hstHxNl9U+mHJDKCk3MxtP01lt1tKLjY8YPA1PIbb+XwgH
Tp1uFuhhSgnfhBhT9GQDkAyoQgVaUCtCPibaWK2P3RZfa/g+lChKkH6vg2Bk1RvsHIt5Nn8a7TdS
8CDI629Z5mHQlgSCWVtLb2iQ99UaNAR9mmWEUwWixapKDF4LhhG2mGfIZ0tdfz5qydUaZ2LdSvM7
a3wPE+J+seU+iBockJ2x2iIKj6ttdYOawTHsOiHZg7feXt3oW1dGfwGhXLV4/PGTBYnTk+JDAyhS
H9TRqJeRqRocyAEyF7KW9yKZalpCC7q1E0L5XY7S7cBelvOLHAxzWjb7ci5dezAIVCsLOErImLev
mnHFHLIh/fTCiQuHRsile4rTx8SPmyAg5Kwzq3HKrta99SRS0a/aK2cr5uzyBFJ483xwYfyPQ5UM
UwWACFe5t0HIrXX8j72kgGwWuYbTHAeD8H5I6CH28vCzz3/qWIR2+dXRh3Zt2hA6X+h6vlJ+1PSc
/RV8xcPodQA3NpYnlup436UmzpTOBFE9RXnKFWok2ugpQI+SGNIp9JPJ0UWGl5KzDeum8FCTT/6R
c15gcysbtFsZN/mR/VVavglZCUYn7oneRsUv7vVLtnnXwTGAd1PI7bv4dsOI51EXOwhA075iJxnS
IqxuxvfuDnjEqZJ/orauu21Vv0P8EcBBp98dFRypOrGdKfmPlu0r6iJGlO1xOIKpRSFu1NL0JiCH
5VxOxa0a2mm7oT/Ljdn5SQ4KLiBmBi25yX+LNt4gG5LL+Bqu8swQ75LXUxuQsJkX5m2QP/gzPkDx
mObhOtTfr8b9Dd9FMYY79D69CBQeJylYro9JdfrtEf59gDTXEUuOcoM1DPJDQSfptZV/gv5StkOl
gPMATT+xHF5ine3GycCAbEgPBCYOoNsXxheFhyTFBd3icVPBBNQ6NnIJEKyJWquJ6rWPtLhfpnWW
921tiZZjLGXaPNILVwaMLu6icDuoIy8l0ks7k0xh1eLeWqhaW1xC78qUoSf07USVIMnNprFTH70O
qtmnEU5wJhtLZnyeRLAH0WkqE+T2S+OyEAXU/CKSGzvw9zo97t4wWzO+GzUivQdwmpSllaUlqUu/
f4/IDOfLlaokgvJKj13m2SlpXwtq2YJ8PSIfFKaWE/f08YioeQw40dkd83RK2ENQ19Xk+9Ld+VU4
/Zta4/B3f2XXxUpQpeZSfJ2SrsunAcTj6RA8cvoAXozD6xP4Sm8dkuhiMsDPBJb1EVDvxYYNckdJ
7PyctVX84d9tfexW0LinGYuDrTYWdfwR675ZZpHEUUG7UQEjkBS6vevqCaIRr0T0eRWqng6H89Kp
Up7vuX7pT4cKS/WgOTEwbZ540Sfe5gWFD20dXvMD9slx7ORGGEjUv95BzDCEtZTIMGz3Undxfy/G
lB6anNMnmPuO44ssJRGSeYjWo9bl19y5a59LclVwaVOpcyW5Z87JHzkskKzrIbVLHCSt/EqhZIAO
iKzN/TIccuu9HJQkM3k1eRi9bgot3P/Yo9qqcuJf57rUnbCbiQz2tRKoHmDZEGAkm8BArHeV4fMe
eJzwLmJXVv1/Z9j+Xl+dFDAuR51rSwfc7IQ31FA4tGb/NMEGvv0iwnmdtQ4Z6lF3FeSyJr5oJsHR
rRqoXsyNDm7zOT88xrA4RNMY7jnQnAUQxD5mEusGDd7KOyAaDd/re9jJav6hYAhoOyt4hb2jnkbJ
BueV71BTW7ScoaL5MqevgqzLVofRu9IgEmcAVjre8TX+GiDPgz8OrJftWJR6IaZe/Mz/eh3wDo0q
dRGg0YkqrZEaYnnVVaqNuMvMqpis0AwNlUsC95JeOuzvrb2YqJwALdkt8d6Am0fJAflxsThyl4+W
C69sNc0L5SoI19v9TZkX6Q/YIw/z+tOrX1E9+kdpUrqtlmtW2PbDI6wdkSry0J++gjYEE0YvE/EE
SeED7r7i3rl+AGlmmP4gd9aaF13SQv4it4sPb2eVavBymipGw0BAlWUV4zZNXZ1n2bkUQOjwSVPX
FJC/RkBCckd1GUgH5bSQqbhoEsXmLy16uFrSy0ic8ft2IBrezq9nLQcPvrPbIsahWfnefBzGoZsm
l2fNhZka1kVO1Cd5dB56ROgGcnrlXr4QZV5ptlNlgVpqQEJgTePCX7y01Yur813/wGI08tRVPsLj
I5stYbeHq8PY5XEybR4yB19N/aeKwad6++PhpOZveuDdKEQs8vIPbSsw5u2sRiKGLI3re6t6hFdF
HZXegag50b+ySpI0pfcmsJHuxNzz2khZ3bGte4TyYaH1+l47DGji9wG4sr1o4jD2PGuH9S1lnxg9
SXTRx+a/BUrBw0w+P2HOgKHsTU7BSSce+Cbr0so0yBDZapHlD6ptWomAjfEBFOOPfrfn8EjtJL+U
jajwDh3GUFOxG5+nJL7lR2anUKc3B06x7NbzC0lZIJu/GWYHj44FFA7aokLtvjbXXKSmeboTciyE
/BeTcaZN75JEsFaS2ktceItw3SSkMR3Oq5uN4yV2iKUp1ryIC6uPGcB/+q9PCoC42I7aQ+4Kw096
QQmpI1Bm1qzHPxTOCavq1IUogM47KzOXe4ccJ5oRmkJACl1a4eTxQRIQS9zcAkhKa8KaqCeulwx7
YyioNHQ44FZvKV4O3yQvtP3vp58A4I/5rXsmOvGx+gQ6W2D1oZ0KGFxAM5FLk6XvaHB1lDEmfrQS
R9dCv5tYRq50MXjKAwt9bAjPLvRc8zmcH8TMJ+IeYxkdgUCQwA+G2SC/tB2bFsDCRJh2ttdAf8u+
QBFGCMsmwJ0Tlrczt1GzTaZ/jXfGpoUg8Vj8SJyLhaO6Ji7TaNkiOfEQgqX2DI/mtO9SB+DfYU0C
MqZK/m+otCBo2MVEuB9P0b0DdmMefW+2xaxHHaHjsotKqb3K7LyyZDceWKHsj+7i7JiC8SZbyJQw
xa10rl0W3pmwsJjAupasahM42uMr/D4sR9+yx6uTZxf37J10RvgHvHbNhz3IPdTlYIxXyn+r6KXQ
pslbsO8ctga1+UP9cUlzl/IwG1VSqHEy89cpG2FOLDtHCwsEssLDT1+5n5KZWPKSF8ftegFXx+I0
RnYCf4brmnUIgJwAnkM+A+Aw9ugA88u/iYhFWLncNvmmMfn6nRjYvaOfYhqL4da9z8j89yPrJ8pR
TPPbvSlkCUFX3ls/rx9/gP8JGD0ixJK++B5PuLGFFu9+2IcwcGEc+/WC2SoEWzlG0kX9r4QfMfnj
GhcQysfNyC38vm4CQUfrnVJYQ5vBeQgBmtJdMG40Mbe+GvxC8rLZ7FitMDHt7bm9jCeh9qL1aUZi
eEJRXgxHNTYhm45zG3/N+ExMV/v9YR4LThZ9/Y8+V/nphoTE/L29meo1ncaI8ETUhRQ0WlX7od7d
Ocq12jaoWskd1c0FcpYuMNoEzEdYprI70dArUvpIt1Lzwv7Fj9yUqsTBIx+FBME/0jHBkLK4MxaP
GO72PkVK34PJHRzlkZKHLacLBs/a1bzGS+Sg2O+oxE+0YmeCG+kVzyjBmLnscdPM5+RhwI7duhEg
Md3bo+Jxmogm6zm0yzTkbxSDDBGHh+boiqz8eErFtnCHt2aglztbOejJDKY+mw0WEHMcEldbAgLf
mYs0sqTtFZhYOToqpEBiuQobYZqsakIxlUl71FDHH1BGDa38gGTeoucDaGrmDsObCprzOodwJcNr
BlVS0418/OVNhtI25BvJTwf3UHazjcQtmFbUHlO6ZwgJHQrAVTgT9EC8otCUwpblZRn4XIHf3BAB
CNrmz6fkVvimZ/BX55cXrmyjOk8pWe6X6Uw4gB3WXWlAhwGvtfo8/Nc/uyJHJe8SGWroNO4J+ixm
/z3mTs1rEkntnOo5nk8WjkxF+d3muVVyWJ7QAgI84v70biXVbSXeVBFveS96FZZwX/Z4nUgmk353
quBiB8nhDZGXhu14vAx9/d2WiXv64wPpeiY7SHmJ2TA+6SRyITPASCh11D0mzBkAirgx4sb3mBjp
JdzFVX5DPlfUb/HyNq6lRXYarp0Hdxi2iTUyeFEBYzLb1lV/VTF8J8jO5oC3YYg1ztCbFmlJJUvD
dtNfiuJi0U/ldDMCVOyIoehIKk1H6Fi8Q5jqbf7XAJEeAJF8iyrUlnSwGRbuq/EM7owmTQbGW1eN
Dd/oExSGWsoSvwb73E3ZN0SlJxul6T4+j7FkYtbcR/rNDEXoJ8gGNsiHXZlYDo3029wVOUoocheB
0rYHmKvR5+BHyLrNdxMs2qI4pq7N/7rA2BOmfh8icgSdVKPZ6It61dIH35KjGW0SkiCI2Zhm+Utc
bHVDB7wS5QHZcYymjnF0XKL1NU0a9njYhN7BHL3l9LpImuyAAvp9lySC80yO4Rpu9xhN9sKSHNge
KRqd+Yx4PtFbrexjbsOyX024UbmdhupMztArcyAQfaLW3xKDdJtodH9fH0SqdIqVnwWQ0xLVMUpV
ASdQccIPum5zp7h3qMFXw0kpE2JZk80/7O0dtEJvIEon5nn/nGEnT/fbz4Rid3ORNs2cLwnwqo+x
xkQwwb7BO8t0Z7nHNDn5zJn6pP7rhNC1QRAuUabe9MJN11stYaIxulKRn9HCReTrHkqaR6BQ/DPC
wsV8MGCX3XS+0ln97P1vjExcIBbSpuHqMcYhU/ekhX+S9aykYpUuRkjjeXcCkedpW4suJaam/JOh
MSB8RURmMjg5u+xc8BwpMNJQTexzaG8QAYIPS4c35R0Ya5Xh0hnGq985NOvtgnJ4hkuZQvZEKfhC
rGXpXGQ8MW1FKIZ7C3Lp/CuCwjKUpmJQE9+G7CNZ+NgqLBcw+JzzoIWBVSjHnFVVPBaaenG9QlfO
83UIWkLJaVVDcW5ZCxx1ThTtn6pSGnzhK7D6/glVK/ZbIMmdmAWgxSonALB3Tv24owg6dpAM5NWT
0oK4e0V7p7ZQlE/8Kvuh/RB5ThjcA/OxzNyMIK0HAJuEr8fd5DeUKZMPpI0dVxTm6qDSLTzNaWCS
HRoau2HCe3bkhinuTsB/2ttK22BSLFLuWO7Q1LNryAx/3YxNjFLPr1S8dVFONPsNj9QV6H/hzhcn
Hq/7CtCliRK+08zp6Wn9kkA04f1pZoQBXYzHAQIPeXjGSKAfl/9dG+ARRLnMsDX6Ohj+zB4reZMi
Cwg1XAMayvEyO6gSLM2cQ5H70gDzY4p7feQkQWx5BRiW0T3dXiYZqeGqO/0xJ2JTJBspu/Jw7n9h
XpkEkoQLgxC2//i/s3Qt73sk6liS5C/1Ya3L3X0t4n+RIT3uAk/ILAPrL2qE5JJ/rD8rYagw8BQn
pgMLFcew3WIN+VsmC8J87NqxgA6Hr1mvyvogls8HS9KDHWS1NZhJPM24NhT3dZWkX9UtQZZ4IGP8
yIz67TiwldYGPVGmb4lTqpROqFgw44Ch95DZ6dh58lUEB4xA57PXjj3YMYDpAIjdXtcL250FIVvS
X+x8KzODKw/xwGz8irFNQPZ9e+iUw55r05ZZYFrj3ORI1S/VG9/AINP3ZZdgbjlJPwZnc9neeNBr
QRisxnaJm1s1IFgTzGOXPyfH7sfnEIoEFh2t0SApkqUbamOCuwnH2l6qaSYOhgERPlNNbZzpSUzB
JT6/8YQSyM72JJC8mMTCBcUH94PNso3+6IB6cgFhsKAgdr+YDw5ajaCFmyeMLK32NvwX+ZozEFMY
cdAQ8f3U+xu/rkvs8h3UFEh9atZ8sbBSt6GUcyTLigQe0zVjKp/p/R2OvHSvWvzEnhCltXvxKyNe
FyGEL/OrXgePto/qGBhwHqFDfpYXIaAHoIOcImpLSpDeOdyIByCoqClVVvjMR1LNFzjPqQ/6DxYh
hUlIEQaP0eBwqeiTgVgjp3yyiH+lzOR44WKXZH3+M/FT+6y1VvDi/bj3+PrYNW26bvDvzXGm9TQu
bN6xBdHc4EJabnCENM1B9gKnG5qDxvEicnyWdXaJQ62MNOw6wKhAaLSaybENqRZA6BuMHaqPj6sO
UIFuY6WWgydLtoCMbdDSNLZ++4W6CUfE9N3PdXL5CLuDx7kWX4rUekYCQ3rNPyZ8HQ4/QOsnvezh
aDFf33v8M6k5ZhfWhbBYgds8nx2oHmn+F0wk+v6/O48ZXbXvRY8uXGsRhqpfIhOqYBiivcDGk7uz
vGsyPYa/F0jYAlX6mHW2AnZvCm2M/7asZ/R51MlXduzp50D0oqqEvoRKl/VvyojR5ZetGaGIcyMf
bldnLzUOyS78oWeVC/Yov2gHklKo57mk4HunNzO2XFY91GflN/YGFbHoNlnT2T+UykLYpw6vffgH
f8/OZmPToslsEbF3govHnsnFOkB0kdKEB7NHs6rt7uSxbK/LpAfIX0vnnc9hqzP2APcsALkBZU6t
PSrottXac7i1fwpq2aZ7QFJOMHKwykq+HTUcSMgf0D6vcxoKmbNvczpQCUEk+6YCCLT7XDZUIU+c
oGL+O/KETR4tenIm1ChTkKMnHu6Smoa4Zc+0jWdqPXfSLHvvjKq2EfTX2Lq37YM6D4warlKXRZcj
QtQK+sXLge2pYCGrX2wLDCsGFzfEqiykxFvzpXqSPF/Lr1YddlbmEk0SQvMpmHDoFZMye/wcylbN
CspyWqomil+bvfBqdoQKO1ap108qEPLfSaGtfI8JQFR55GsEmvcEGHiI17F9ELIrYu4BO9oKPWi6
PVTEYVqpMx9KGLyHykWya6TID5WwYCs10JlaXKWCv5KA8F/q7qpGkJFpUojSuHAMBlXC5VHAd8Ad
ZZP/SKjXmsURMoiG8Av/SguxEcdfrd5fB9D1foB3o3VtT68yqv9AT8ONw5/FNwDhwUM4c3VKfY+G
AywrM0Rmt5vK/2adSs27Y/GujKf4Bbb++gWqLwLh4xFcxakTm0+OHnU7z5lvarmCOSIgOMum5ypd
Ib5rMphAjF3Mr/vPiDIBuhiBMB50gRXpdHl2rK4XYIQYHsPJQNOJ8Js2IRIPEsJCbB2Zv6r/8OIt
Dv+4enpzH/jUg9IyVWYWKk/eUhEC9/qBNCtzlcIEwzWR1fIhLI06e4ibK16/qFk7HkpaZ0Nx1M66
wWjRq7rG8aM2R7gP9VTVBtJ9wGIooYG3m9eOcYWYX5ErIoT//VKLLD1ubVKvODfJX/a6hyu42JVT
YSJeoLlPqBXnR6PRuA29ai97At8pBMRCCRrdj/0wy22Ow2+8i6s84D4bl7JQWkDz/uZ8tU+dKb5I
NfoBsZMTgJa/NMG5nu6K7A/AnuFc9sFxHJGRSEtaCGGOOZPQqsR3wk/iOr8VgczrZcyKXq2whdtI
rxjdpglazGaJs1iKvZu1naFtGGdIbNZS1goDsNTyDLb89VQruforteiWJWaE8kZytut5F0fief8T
hGoQykryxecXQfOFCn/XXhlqA/XzQLZMtk6P2Qt14burmV3evgbWacZdYd1X0BG1SXdqDwkQJXzW
TwWwr+uArVfR10+KjpORTRPUypksow+jxmHtQAnevYfREvr6K4UcMmciadMApJwY9xxAb3c3RChJ
4hm03OO4YtG8NYsTYCucTnULaO0Epmy+t6ZfjKSJBa4ISNv5mQ3G7tWI2+YR/Vwkmnlhc/wTXJzG
xau7y6lHFFlSUZnra786EO+PZJliK75e2iM5LQRinA3udIvuxyBhmj3vdQk3b/CbJwQISoYkI7E4
rKVASG/ukehtF7bDl+8NO5/Df/rJjzG8WPRmkxGvuDg2dyRB0trXi6h4e4dGl9H1rePW7GJ6lgH9
zFHbtG9jTKNZt9tCgC5Xbw3pY+sb9rI5ljaO9p0TFCczgXlxvl7fnj2TLygp8bnWyNn0s9cmnXqt
9wHofs8LKV4kQcbFLkwNC0SRllA9AUJ45R9GrsGsygwYuep0gTAvuBZIIsqSLVaDp/sGzIt9QjlM
V+Mt3ZDLqZMNRcypf4gVisW4+8pHh14SvqIWUhOze1bO/NED4zrvWc8h/a60r38JMjtxpUnEjCj6
VoSQX63Wx+1P15j9KdnM4PMOjfUpo90CcOJHZ8Rl4EA3ERoBvRcNu785M4TJguKHKcOrnaMN0ueT
66R5PbcYWdz+ZLbKw/QxZRGKWygQGAtRQDXuKm+Clu6grwVtwpxhWAjE0X+JPWGIImwDcl7YKqYT
Go+Jsoz1SGdf1rQ3rQEcU3eYPCPe8KROFV1x2bSsH8UkB1/KEXUeG3UW7/xWpCbUf0Uu+uJLwTcM
nXND+pIV8rQdpXg+hKi5fR62z2s4vGPiD8ob3TpBUoiENLZ0iM7+HycX6pbklYeh53wxw9WhDn+U
17VbALCIEYM04bKx3piI8rCtYoBKbh14b+vTRdcjb7TCxY/QoDOQD+Msj2VtvNFJ6YrwAJO9Tz7m
mFHKSsGqCSNOzwWUYDLWqpp2Buaf1sOFym6Z1uYfS6ha7F8Ruo+WOIdfV/SVYbZbKN6SI+sq1ibC
V+IrvsnhprWTbMcAm9o4IdODaogpEQTT8dSQHvpQWGKv9gQGaaS1zPCkV/g9OjDjs/lVBwEkiZ9j
8U2fVXN+TliSPQU13Uq+TRul5hha8vWV1mEOfGeYNNh1WXur4AU/CcYnXG12Ekt4DP1ENZei4D4I
oNvXkX2Hmiphr+M/pjx/m/lrpLSp8ewrmw8oFg8dP1bHpMQk8Gj3meQLu1FpYf6rOsqw7tokqahe
AfNSTXzARwOAU9tBIqM9GdZcAOTDdo4bRNg+dItBv2v4uduY7hu201gqxJPu7KG84jgk7o9t4ZLX
MyJS50NmZ0rXFXu6iwE4wqwpTRzO8rEfJRQq5POVxBoeiDg94Iu05UNGVY/5p5hSxVt2jnAHW/sv
aiXUSdp3nix/wq31geyXaMC3giLTCBEd2ssKBhU1Q6bduL0RHMYLMEpQ391Ufx2SCrISLXWdpAgO
U5hrxsTH8PvRA88H3FZSnnEoBogFV06YV4y1SiqetASbi3XZRq/khYhf+o78mPmDMUyBrZBdl/ym
zISkmFjHq+3j6YBWSRO+xCW++fDBZE03+5Tstx5JjOVlI1Y0peGlvgxu+8OiwDl7T37/uo3lHbvf
u9dNboHhXRNGCha0lxQvYreEz31bmblQ/pG9o1Bf0ZrUoB3DEH8OfSeCFXu3f2BGgHpFT37MV/3J
E1M/a9t5p0NTc98lnbkbQQfvggXeLcGL1O20rV+qmL82EDDmB1OBhTG/OepieeOySVnlaK4hQ8DF
pTRwMfwv/GvtBPOZpX7WhjdxUL0DTidvgvznaHPhFvM2otbOzEfUojJx+0o6C+lj2xEwOH5glvTi
xtb5Ny7kYtZ/T0xX9NrmQ2n2BadaT8gGB+QKiSkzXwBh3uXF09FbbjUEPvbOF2duwQURroRUrXl7
ZnVWkqtx2llvluWfNZW7x/hnW10kGaliEOI1Cd+IECoIX4ChIjmW6f0tNK+UzliUpQq02JRS8yCA
Gd+lOoQZSsoRKKyRhLzgQ4sk9KEs4DWd0qs0d5DSIWzfxfr3uksw4TF7Jjcq57lgXxqXjL74wKU+
GlkxYEFj5Mb70dOHqXUS+CKQJuItUlibGg+iFLA36e41HZpdltYNLhFbLBJnBSecn55bWEqq4glo
aJLaTOaIUwS3YvrW5wzpG2K2sKQINe0bk+ASTESqpBEFW2uEHo3Z1ex5BCxIeWBO8/CGeDKYNpKI
kA8uVSVJPzjsbUkHQxbVfyEjbTlpL63at/fmB7EwKKZbuBDA4bpgChZsGj6mFMdZRE4vwDEbO6CU
/iqDnXdnysX20SBq/HqLx8JVHT+EshzZUS7+vGlQsIHTzSaJlFdsa4zRiqaRzIxrqc7w+zcBrcEa
QSKNGmC/2nsHjuE0j6TsNgdzdOPuu2FIatzg5dzDzaw6PydrEMebC+ERR1Tvcs1rt6QJyZJcpAOw
4CTfQgYfLy90HSS2w4ajn6O9xJAotWsD2f3ewCLoqAuV9yokXaRrNhKbSqwvP0dtij9ub7Rwu1+9
gqwyoSe1c/KCbAjODO1FrMYZa8WpBT82FKc7zZxsiQJUvE4Nt2iCjT/Ge/FOsa81VcxZVbcXVKVl
g9KTJ+W1YhBitdxJSgCbBf9Z7RE1+POQkbPcKOvbatn+clCau1kSpVCVdRA0YbqPF7Gmf3n+/mME
AvSCvId2IMC21ybC7xyYCvI0cLgmutvloPbzzIPKAr2cMWp5GqeMrgwVj4jpvlOa9qJO0YGy1NNv
CuSi9jl4JvNnVV8Qyz+rGwNLKu3tFU9gNEElerk4peVA/udNrC0v2EVie4VktU3FlWwim5y1UGx5
owFCFJ0+74X8NkqpOLeE51euX0+s4wqOBrJxUBfjGZhHX09M6+6cvFlzAn9u9shm42yzPgzGtXgP
W67ReiYPbNwe0bBi5YrHBQv+EvaeiXYWW8dSH2jhV4etou4Hw/DaE+tH2clXt0m19Wwv+AULoMwL
wxfs+yQDPsQONIUA77XRzk+vl/tIjZ3GTLU9B8goPq8f7asoZAn4hFlgIURYr350WBZAkL3M8Fgy
cvqcSW2yu3Y0wjaBw8EjB2TCs6lVIK3Mb3FddHi9ViucU+xvQR7SiwgHw59ZACpCxgOnwasa+wFH
A1ZqVJ0maiLSZn6A9Kqz0HGtLafTABOfeKGX22qvPo6D/BJtj+1ReboazNO4bbfi8v+VB8nyafKg
x0yC2sAdPTa3ynyWzrzwMSFdhCgjmEwMFhNNrI12DCQdqRW816TgBeCl5HWH/i6bUhgXAKEpv0ZY
FNuLBd8pYsjw/Z4hTpOrR6xehiy0+pW+Lyf0YwSOkwo0hY1gDtCstp6y3SEh5/jkHUB/+apOzxub
Ezi6Ktq0IlayUFhZVBElppLo/0eB4uE5UOUL0N1TlPeTK+FZzLTf5bmFCIP2VMjAbqVydmvwP2JK
WV3mk5YXIGzTSYzeNi+sbTPVx2oWEvo0m9IrHFuDORRl1c7CjhdWulFfC6YoFpEEPbxHA2bk0RyQ
QyLGRH7RQaz3F/4GPDnpmbyBAFdV5ZR0C/9d7iDXfyszTlFj4Hufc7LYKUedm20GqQe3KnDyoeN3
cDoa7vuGm22n+aMjNYTG4o2AgT6wM+sWk9Qhmp+5I6iiIK6NJwcBhQ+ykGiAxnG3foFQop8QwW8O
HXiGethsDQEDRpKtsk+E6EZcmm6eha8w7qtcnjboOuO/1Lg4ks1B5Sy0fMczaoCFHUPF89O/JBtG
XhaUX1ULP/GYVonhTBBDiPcVtsRpvAXnSk4ENNYrCLi4/aim+YHxe9phfW+2mKayyBJBPO+7H5Ch
K90ukBhNaBkoKUxYIuhfCs9gelloO0IyXIpeB7z8YjIRDygW+i3v83wynihqQ4Bk8Y8grqpZjhBt
XyJGBklrtYcB7Try7tU13u7eSGtFnW6HVX/hyIcpVlkkX1A+OAH23Od47hBAzACPC2yazHCkVSwc
BqGxW7UiQpHfgy9zVUaZIDfNp07pKlRmH3IzMeMT9nuWi6HqTmHqgfGKgFxyunH8pfUIAtWEB/mU
NY38uXb9uPn7G7ICeVe9uAsGE9CRt/eQMUpVTmBDZAfi2r1ZA9aHHlSwp+MopAfwqQRgzn8Kk8NN
bd1+8la2oie75thmunAZcrGQMoq+SuHIzpAUhr3AUtOVqpJxYyl2WZ6CSF7qOxgNNOXD7DHFvtBL
RWYQw7SNAOffEi6e0XPPOLnnii+vHXesG5wba4T4r/NQMf/fkcviv6gMU05sRk91H8h/I5B4L4xS
YvJNfa+sceatPSCNb+HHlFLO7z3BDh6WrYInkhGoB1yaYPEGnNQHHgYhsCy7oq1cOHLfc42G2vCy
oa0/KueVQcg94fA8pXwfmwZx3Tikpp7F5Gt63tO4qdW5pUXq9h0J1+LH/fN8YcMkP1gwWYZhTaQe
ycdFVOEvd4ZxLiPbu/LT/4b7ATPg2B8zhtE7X1S88aSfLzdEEGtrCtpUDnpbswIa88xu+shCKsqQ
brvd30Qb/JKBHsUghOIcBS37EqQCZah5GpsJIbM7vS/PeMlwsl6KE4k0+t/yTUFgmMCarY1tKstS
9r72P6i4rsU4ZsVS/Mjtk4Gk1gEMXF/T4kj6bgYJvuVDNGBkz8YQTb9skGQ8OtrC3mIWh/dIFRW3
YlaqRyP2uvpuJ635jpKt2uQpgNvOUnQwlkwXvSog94yF09rjpSS8wNE9dUGXHzHREM71APTIz3e9
zlDtuGclVqe1+3PZfXPVD4f8e2uaCIDJk1m+0PohQr6jF0tWyLsFcaoqygAXGIL+85XHiHDQ2J6B
EPlmbG0rEfueS4eMvtBbDPAZzJXCwBaqIMMRHLdriuXeP6NpDEhVX+yL+tXwaF0wyTkPWoNQUTzP
+M0jG0hVXwGultruHc2rpV1Byy9g+LrWR6ku3jxaViIGX+HIKrwljuXrqtlqVQD3I3xDeNg9urAh
D2B1cm4E5iR9LRcYiDw87LE2RlqQpF62uWhTu4TonMai+einy+HwGGnItpSZKMFa+LJpaYwUDObd
Qszm7h1nxvz7noJSYb8G3Qh+b11593XDkspFsXlxqaFxc38zS5evJAno5Ca0WtFeTY5ocTN+aayF
fAkybLBNMycJ+Dd7B+20BF+tCvrTq0pzI8EkGLJh9D9U/evTGLkVWGCkuUex19oR6pA4bjVWIWKZ
jevTCzc22zYdx4LFOT/C+KYL/Z964X6jq4rcoAtvhHNS4fmBlrBWVOeJacHbKort3oqcit3F8+Dz
4v9FnEA2qbyskQFwJfwec434lGbq6dEbvt3VqTlwBFPz/Ka09rSaGFwtVMl0S/2911UIrQF5EDWB
ckR8ZovDlrU1mrY0wGU8XzHPYccB0Ne6KCu4fMVFYYzzMEoZPziAxRos3mj7uO/26RBWND0GGd+Q
C8LusCCSGEtZIomscdeDdh2EOeLX0+Cpe9J0k+vHJZRQ6Uba55GGhu2ScX+WVeE1n0Q46PN+etez
pmwGE8pAAPwvpD36NfzpL54n7yoimP4PydcYIk4JBSCK+7gmtW10YBUrER2S1ioDw/ovAg9McuAj
o259PMCxClw7cNmAUeiUudlMcAfxI0DWFjJDXFnFDvHfXX+lggPSl6pi63owGBmX/CdNLT8H/xwZ
cgBeAIZb2hXsyuWyib8m0b9GquZ6CVMRClmYLtxtrVIZxwa7fBEjdYUHZ8lWjdVA8ZIXaRDR3lqr
KvYlKFo8e8szJJh0I/Fz5TJKKV0Gn22txV0fzo/2lYzCwYTwhheyDUtIBLLd8X56DgsMSs+mOXau
8/eAtcHPIps07ZEWs2UfauDsV3H2K1DcnfFrdjB3Vxfx3XKRzaEfWkY18w3uXV6XqO3Ay6Trn9Dc
dB5k+qoK9BY/7P5PwotUGP7nawqu6gbzP601TJaUQaTQs8KiKubu5WL+wVKomRvMrH6LhEhgp5Pb
eV9YRFEO4xSrrivUYBUYr8ePX0dRGfjD/H+pFWg9vJISFNembc18d1VYRVVvt31rxVO5jToe9KQU
+DbYUf/+UsDGUQ5ZwZIHIC48TAhwZr8oK4VUUhcmKTZdxv6QPNFGUmkvN6MG2CMbsyOZd0tmwwA9
l6t876CUOYwsqamO8ZeZ1gyRgC61gHnNfSiPg+TMhSKHZw7TXWbh9gGFx7MOdr206504T/ehqw7b
djzEzSaZB4K9UWh8xluWDXLDIMte4Fn+toTdbR/m5Xnl4txbgcRkyE9BjL+rn+EsInIkQaykAhaN
lMHELOQJNStthhnKlID3I16eU1KtGAurkMF4t9ijX3BbfStTa5bIBjkxM0RuWw4OzaG/+dARtrtG
z2f5JX8Ozpf1/zgwnHmSdf5QUpr0lErBaCAv6Fi3wtU/6m2tO+a0ZUr3hHjCHELE4SuL8kwNlmUY
gF6LCyvDlqLCxCbJNMi09mTvkxOvAD/WF8f0jRgQDDasUfojxsGPBhAKcoZb0Yds/1ld+UyIM1KU
kSAOPKWXgHYooRlmFiiVvNwuB/BZCcC+vafJYbSd+7qLUdvbg5n9awtEkUTOw/+jPl1sfUZ6SJfR
H2IlealNkSvNovVZxXWC6Tqj0vMJRh8sZJTgkDOZtdpqbeHeceoNXf/3rFoZpxsvBRhKxK2YK6Uu
NnIc4PFc5BDIzYJk9ULoGU3k2vkmdSNwNSMtJ+rak+iubOpvb6srM72tP3ntfAXXNYJt5tvf9iEa
fnTZjJEIuDg5amwMq9d4grSEFye/WqElW4BhOjuJZ8RQqfrYa1ObJpkh9bi77Fy6EepDmTNi/Qkl
s9BuOTzms5jiye5fRL3CtwbkD9zq1CreR3EJE8TFwEdvzX5yzHdu38nOkiYEBHkgPi3fli7SXEMt
+OPE1OAZczKIuAPwervG0nTt4igRXLQnahGsK+jRHsRef6Rt9zeopNmXBXOYbpBUDlfy6JJE/7qg
3qtKiUWnHT/LVasHFQY6MsKDCCDetUCggK1XiHnJ6OC4MQ8UGgIjN6QlCi9Od3Y5VviCc1xdIoZo
GSwyQUWk6oMD5SM7ddB67JTDYCKlekWwjsCuoT2b4Dsz3O9QQZJoH7Jz35g21/ifOz7T6Plxp2BD
UBwPh36UweKXcyD46CVi9Umeqt04xPb+Ue/Q6Q/iuWqTdWBQritpmVBjVhcNC0xD0wV8OAnvb9Bi
lrT6ecblQRIulkjC1oGIwFTg3Y+JIK42v78eYglVR32gGRd1QJgf73Ysz91B2lCu6mksQ06HkDql
8tQ0tcIu15NvxjtRO8128GtNUtL9tBz0bc+KBLGAZk/j/DPOo36WeEe6s/ZeMGW/LuAQur80Bws0
rxrugPWDgISSO/Ko0MOezX0gYl8Fx34D/b/QwywDItRGD749XnAt8yM8QFV9Ih5/jlbLbZNAuy1E
DAlAhQen9P/qMd35Lv2rKUGYm41cOqxGxVzatZICQ4XpPA/RJPCHrYr+qU/2SoU1RMoZKCoX277U
V9Yr/zATnh0KvAwtyT7INqFkfP+1WIloEvivVhpjmpk3WBfdpJpVQ7YlcGYNgn397QgRmqsBtkYj
/4md7RRlHHKhDdfh87RteKiItwUEzZuGurRtjdzrcXodkDKea4kR5qV2sqcD1iD0j81U3lR5/Jwz
gWS0/59yJ3aLbGNKyj2DTIzxcUqnsfYDU/wrewI/i7W0Tqk5vhx1RDSGAFMh62KmoY0jJILz/k6o
cql/v8fdN3Vpmbf2i6zCEQYBRYNUPZHjTkeHoBgDBJyFfOo1PprfXpWj4WNCROYgJAI/0UWzNTUw
SMbMJrqRICe2ZE2rdF1CMoDFvPOEwxdc1eT05dZoDwBUHhTnSi945az0VO+lxbgoqbyRcM0Ih9Ny
aYvMHRhGGbNAFEfFKz6+DlkOJMCqVLeqP6b0jx3luc1jbk31GNv70pSn/1Epjet0Fcl9N+8GeLcA
nc1PzsG5iKfbQ7XOz5ff7AjMxyLI1ehypISbDMdvl7pAVYKxezL9QotKQiJ99cW1s7KoztPkUl43
ssCbjrMZlo+VfDgRrO3fK9fbg+ASKDmE9mqQNC2HQEGAGx3tRocvmpOY4XJDfFuUSET4el8TCvzv
Wa1zJSyReGp9Gpyn2Gjzd2Jg0g/yFeUl9iXFKXg4Ol/oXTiysa7SV/3bAxjXMmqVIuo0p4e5N42X
9r8x74my01XBeBJS/0O+xfU2k9ItAHAwpZ9bo1JUXp9ywywLil6XH0d+Iddj2lplirS5hk0HDQOz
C1IZJsWSdP6hb+0Uw//puOLn9IpsZLej00LyCAcIIk6h5pPGw0YURgp3DI9TW2UgbqICUknOLVwZ
6+y+HhiYaYYJF64mbOxpKmFEOh19i3ii35tVBUJcIZFVdeAZfccZ+q8OUALVVld0Iba/vmtYW4Up
UveUXOAolSJJLsAxFp/3EXGczLI5XhqND7CYso8RBHTteOKmcCCnfa8pLgBB71eUMM5I0/00SsBP
2uRlQ06ZDXlGKbut/6lGpAVGb0UgZep68XOofS9YSDwrkRwgKzWlXWWLf3ljASCDjdyBJ27X0tNM
XN7UhIMQMvd/PNTjXH7u+OPy6aD6myKDadRLrLqK6NEfrGaufS3dz377z6wlJf7YO5mP0DlQIq87
RPSJCznE2W5LSZ2nsT6cwM6kK7p/d8e91dHrfK/3+kPlpBDv24th3haChUFpb8OzxgiotwG9ZFPv
2szRzxeZ/p8qi83jg+ctYMYphd2cMQtpZcoNisHxnE+Q48mLQaZLzWA0MHJcP1aikZxREn8ENqfn
bu5v20EiE5Ij8OLfP7PS8gCSc5vodB1ogmHqb0JjdhB4K86ReDp4IOocC9LXJi3YRqm/N//gm6dd
q3Buhs0+7gS6STHn33xd0/ft5ybnkTZTmlRIISBn6kjycu6/BH3xnSWCG3xaTN8em1ENM8ffk7NS
a5Cr1In/EsPVytdf+sFbvWHOweNwp5w+oEypQ/wik76xy44uOlgKj/yW3iMbFYvJHj/P7T89eCKI
OeAsN5mNDXYys17Ob94bbsQmt4mgw2TY/RPAmR5DPVGrbT7NWKjbgGqCCL8B+JwHKhkzWdsZk3w9
ubs9PnHSesFL7QtctKOWF4kDh7mjeE+QDdWSFQ4UyYtbPef66H5fYPBPaIXi/sHYDYk0uAsIIzJh
MpDtwBBiSeatH6fUD6LZ5zJeH0CLx+8Dtj1un8TWR9IrHgS2VO8XwFmV8/xtyNDIn1rNY6UmFVOR
JSNv2xDh8v6sqPl1svGTsH8hNdMXD4Q2JS/CSugaylah9p34wI84A8BN5TWkznmCSc36+GM7CL+T
QKzUWoSLiLkWgUFStFfdeI0KXZcvMWvvarRpRuZyVAOc8/d1f+k3MDOgKDJBz2NF3pHXltLQLLhO
mibCFy9euPzwPRV2UJvm/8GA959KFOGlyc9pZRMXORhvkujR8bG2uGPferSWM2mPdfbCYLCHVgyt
kL6fY5xxFRMDyFQWQhGEuta+bjZZ9GJ4+pNLbl8332kQlXIUmB3nYDP928a7pSUSDbHgblJKqrMp
Mw4lMUckws2kAcw7Bbe4iEHfSeGzNI6+SIOEUfXR6x8q9lh876B1bfZ65AfPkyVAgG+PcnbtAczS
tSRBkjJKxn/9hvZL4K/O05FiPYyFHzQqtrGlLBYQPEkjVLDipTfOetKzvB3CeJDqttem6pncdtJZ
c+6em6/dOnTynvVbKKAW0Hg/0veQLTM+c8vqnCea5aC3e2c9mxOVR88EQuB0SrIrST4jiCydvW4w
p+5jBcXRYVtksF5pVcRnwyl/lxa8NyCpGcg7O5C4RwNfMMHjZizVcXHhBluzId8QO6RmFGlHzsGU
nRZBlTecyMaWJntsUt6NG9KHFWHgc6UETuFvTxv6OuHDPvEjeCHC68JZSRWTsVDoATfTLzkP6E/G
SbxflRxMpnejUcQiZz8R7ULknMzLkK+JZXRyRAAkXBuKz1jshx4B/GTrpq+mCcmYM62rAf/uizb+
9yPvtnSbXikT7kOxfDNvjMs43vUEbcEP7dzUpCeU/BiIC2xihqrXsw+PHfCKvXTofKWRRo4M2KSG
R+go2UzpUlPJiyHh1XviPJbRLwcmYDxwVOrQ0wcgnSHIs6/dx7aHoB792duooFlDj3TriYmRLnk+
RFg/HgRtwQMIv5iMuPR3bsyfMTd+e4IXyr7S9eNvJ2PWuarVWNd3a255djMQKVnZuBYAi4UFeRK4
Xki7PY7VIqfH/S54B6xdXINFzKtw7EE6HBbUhXAF2jAlmHvVPiFxWw6JuXZ5gqfMTWPrPZAOsjHB
/rPMFpQriW+i4wfcywC6WR+wuWJT1vxybvL9gI3ZTBRos3EsnUloQ5rYyELQVBsD2wRB+YdP2n93
UC090w6T1qHXIRA5PXtJPeFDWWhVjl+etVIsaGpjMnug4g0pKjDghLgeWaUkzYWCnWZ6dPobv6lO
uQAjtQedCZ2jcUeq6zdM7ufNZ2xfV+ugAPzteVq5FtgvcqKY78stqeEnnJgrRSLSdXW9UUl6xNjn
8eutSeecYaFLvJrQEeQdDMgG0A4oSWRNCTAKf0yodHttwNEbbLp2xwYWV7AMxD3xTQp9Hl0nxL44
Eb7wxvSmBqcwsdVQHDK+y0wQgjGjRCMuOloROAi7TIQajJRI/gI1pTiZ7OHcElrGiy5M80BKRUYg
wuq55MfZgVUGXivZRN7Kon83R2n5buj+iCejWlg7Jv71dLtikonQpNmwS45d2KjvYFGHjIAuzqrM
McOD6V88XVmO1suT7d47dAPUTDvwIl5ScMsE+rpoIy5QSKNn8HRw9rXz8FebDWP0q2VRB3ZZGpmn
EMUWYWyPxanvxarjoO+nCCv7Hg3gM7U7Vqaasl6RiKNCHtQSTRg7cKTcZ4jOJETK4bVKV5WLu9rj
W7/2x1USwMWQDxuEo7b8psjy+DW86RriXADKsv0pC34K/in5VTTcAm+PRkUfu7ucdUufLz7iUvew
9MHIgwe+ys8R6QbiJalOV+VGfeiFm3zTuH32wfmBR19qvhXOUGBCMERMki/nA71GCgOvwtom6HrQ
HnboyMwA49C29Ui7LMyDglIEcUosvkCInwnZEwAr+8SnN02D16JcsjpH8rTQalUuAIvTz4iMrEXy
wD/0cm2wwFBvYLa2H3bn7eB4Z6fI65h1kgeuS1wh3VR/I/7TWESo45kr9uGYadEvOw9q2YCPoGd6
ORiMIM5emBcMorq4Lhcfg6BmHOKAGp6zoWhZdMJybrulMFGopRSuQ15I11JVgF/v/R5c9Y2IgZi6
xtY1il+x/bTr/piHs5oZjUAVsLf3n9mCcxV2TM/3iHQeQ7lU1GKTs2mCo5jtBzk5ojssjtybx0uH
XYVaq21W+5kps/1IMw/on4Vn16BkEhkim1KTTrdzJNniHkz/7f5tRQ0Kv2Ya8VjrvoFYE1MoPVqY
zv5H2Nkkf/JB3616C8O3FG5HQmTo51XN/bnH8en5bCdJ5IReKLngfH8BgO7r30TPLRZpKpE/uH3f
/QB65rRRi6B7kAcFSE8JORt7Mxjihv4zm/hst1NL3M9MyRGhmXVDDtelRqkrDtfeIit3Ol+Rn2Ni
ZSCeoKk2v/JD/4YfXDIy1Tufwb/TExjGgRGywDI1IX4M3kA2JcTBtVEG9I3LxeUIWWSOpLmNh2si
cxHA5kgt/enucvpJaP5spQM81mmH5YEKgx3AsTdkJYdADwEvH84mWBr10cP983+A58FUznSKGz3q
IKNu+ysotwKXAXvxZvWjhjBiTRbZWR/ruFJILb65I9Zi84Y3aKKDD0girRU+pSajd38W1flcZjnQ
2AhC62OsbfMrDnmgQPQdXm5iRemojNJxXjOT2fNI51rvlcI8QCTmxzQD4h2NN4LbatBgcrJImyql
CCaWitTMAgKN7oFaOW22ZTwVHaDXPtB0QybUhwcgOYu+PR+gQ0cberZR2omxMw6nagrQvhWLPU4f
kEbQP0PhIezMtXlVH8JpP069TYUz9Wst+BcUynIGUr6UufFfhcYtQZEJa855+xV3hcbhnnHHq2OQ
dWGNunPV6kJ2wb7N6D3DUTX4smE/n1VgXWPl5dFXEM0/dyfcOZAHPczobBujvySFHMNWNDcjwXGQ
gFdME65A4r8SM5o9ATAUisW1fza1jgz9OXWEFRqvHGF7Fol9HkyXCMDR0W3LbhRCZHrwjkbs2cUb
3p6AKYgEVO+7sn1l+K755LhG433PqIoCreFrXjZ7wx2qS+EIsF/ZfS7wmAXIsIuKqR2QCz7xHpOH
MoSKQojyuQVuoLNKnsTXgOIJ0e6doBisFfkOGaonHLWcUPgmhh5k4MvI0QMQ23iRJfnWFIiA1x6n
MzuVSN7LamLh+ml8SCw/DDCcuDCAhlhmURtUX4/itWakpnD6C34rOFIRbpkvk27vsyV8Vk39bLB9
E0dUZ0PRKfyV817w6yDxWZ0JMctSscAxTDnMfcdOGPra4+zauO80jJznzWqsGVAcS55/bhpJLDr1
0+PX8bjTc/GS+3+ruc4YPyjgzkTjYf8IegDL7YSsu7vX97B/hohm4/VTJdfQQIbkG8XDUntmy6Lx
l07LW3Y/RSOhBEQSSFvCwJ1caTgxrBSXpwmlQC8THC93bS+SNjyAr52WeE3im5kA1YfkabOU6DoX
VOmMm7ErnS/cYNc4hxjNc5l0Y64VmxX13qRnZMAZxitOBg8486UPxhZAfsymf3B/H3OkhTKe+U/n
1gv0Ts/g3SbEawVE3fvQ03v32zE+atU2aGiyMDHzLmovgF7fBn8fq8wR3WifxS+F1F0PvdmFRpqd
UB4vqkDrTv0ECkl1mjCaTUNijxPvmwMzyVmimzm7MrCjgIZ1O8pdiEfPaWzf0/QKFyVGA0FnZ6LP
3pwfS+RXMRXOGH4e36EcI+/+2ghOxaSZiB+5kAHC5/Jv5xIIC9Qq5MtemV8y9UDbZUjsjWvvfln1
hx45Jazl7S4eX1NnQIWSiZgsByBKPq738oBAhMH5bl305f7S1jWP5SFICYmDpy22A2sBm9M4MxhO
YY/clDPm3FjIIAEAqT6XI1f7SFTzG9RX/mdlS4d+0ODSZiojyFPsVA4GxLdWhE94gT6csTleZSrQ
9b/3rLKuigQK9oW2Op6dLRlzaKPNy4/Ff/evzceLlAlHYA+V9Iq3rlDwdjvksWpUZhdJcefX0vsf
N2VWipX5qNrCdWqSiKqDxWy8KsZxJ8WQrCdTPa9FWpnRlaA2X3LWjgQB84M49Eu/lfi2LFv6O/tp
icO4ZKnVI21iwrUMAWauPmASr00cKXNjUN9SfomO5k8EgOH9BL/uSsgQadX2SUjcfpCBMcLJvw/D
hrhkYMp+hFbxYVlrlA3pSpvdMx3V1/HgwlqZ0yRjW/pW7FsY8pegdhiR1dmREi0E21gSj17063Pn
o+qMsMRJs2nbvdfeW2KnWjpjOcDjbbA5bqXCuCgz+IgmsqiW8U2CZaCGGJaWF2Lkq4KT/MtFhyKF
nz5Pqbx7U9rWIvKPWRZoQ9FfLR7bJvCWGq43BrUQmT7phYgldnL6Tx5Qfyyyfl1iW4c12kEzlD5v
uMiKEbRdU+tuhCtMRUu4icXp8zaxoO+1JDte6W+TQwfwt1lM+3q7yVj5VURXvu4T8UIja+jWbg72
DoHK7YZJZsnL63dlFZuSW6lVlSbomzWBXQkws/0+G9b1+jiznnzXoaaBLWEqSltjW/FKEFiJknti
peLEbWq9GFIV2lQiZlSaWwz0XXyf80NdBw1J39PiqUgrOYK8xmqjWXSn3M3BOsTK2hBFtaQ7P4z9
akaWgF/vqZliasWDON554FlMvvajgq2cRrvhdc4Ie9r3e5NjZg2P81LnJUlcCSmNrHlzKgLfSzYJ
eykP1FMLDrSMyDjP/pSV5sGPvqyYO3Mgx5F6gx9LM24OTo3PHdQaxxWfjnSckYqOBKavPUh85DDO
hQrawEValmJ6zP1xJE5BpRXilMcxsstSCqnRh6Hr4M46ZFk6KKPq5OuiZdKAkVJSUSbTKs66ylGk
r3LCl6FxL0Zy2RqBxU3/fRciM5zSob2AFUalqUaTaeq0kLykHtUHV0xdSlwjOGXDJbTlExM56EKE
KCsN2cenm9/0WJSY/i33oXVjyKdttYEmkRDUU9boTK6paW5+hbDkaGHyXPxtP1X+q7yuKsFt5x/H
rOENgOm5+fUmpyQkdqTPWs4+IyTEsIiqjlYaoJ4WeRF7LMhsGipbrgWU3FG3yXDHJca7A0IXLP0H
DbmFcjzeWjeWmiUjxe/UFWyHmiqMJV3ne6GW7RFEGF4ZPmJyH3ysktuOXFA0R3lFlkVPJgr26Bko
KNEirPfia9phwGtldipn3p3RenJs9RxpDJ3472ydzU5rFd8BDiaunnYMNgn4peeNHHRuYnSwMHM/
QKyojohT8PFjaJcpLgKwg5nNJHe4qajdf0awUbcTnIB3CvoUSJ3wgpccndS1P7U3IokruWFM+iKv
78QamGz1azt4v1eAw3ofTnWJt09FVYJ5NnWx7tWseU3SR3At8DyQMD5HQSW6rumTI5OgyJGrksR/
uSa6gloaGpkd1VWKq4D9wXCBj8rGXcKdi6JsEis+Fb2dbZXEA4xeYhU/qqDThNa3iEJld9EmP+v1
A2ALfWtAIpIWrhNo3ZoAj6wDHbOMSzcsjI3lE6TXpTg5YE6M8xq+WDXzkEZXb5i/leyDs4ARvnvC
XnwxhoS1SEaD9EC8PZFa4F29S8ADqLiVw/k4rEHUout3S436pXAcxNw6l6iBJfIbpvBmd2W+HCIm
Xz2JMHH8T/NGezBGBG9pYFnjdskacU7WvVEgywU75CKnAbcCAUM26GsvqmwyRruta7e2LiSRfoBj
7kpc4AyQmyvfIHc2qiTU4+Y6NjV7OmO7QDoTynz8iHoG4WtwB8AXxYcKdMYxFDS5oUIPI4qwocOh
oR3ii9z6Jc7prQkUI0rac8HnKnkI1RU+lDglofe3a/IeRA5eJ3XKjkT4Bcr49NPHN0N9dj/i0EU1
m9jVW95RTLLd+hIbLhIkyfjcmqN3q6yUlxW0wdrj0w1Tl9kmEfKNVMi5/PG+BM37ekftgJjhrZqk
gXS9Xr4XIva/jmSovf7R/rcX4wTkgF4x9haByPVfPiWu9Kt5r/XYFwWFxZwxuNBMzAOBfphHd916
uQxNZ9deCAGFVpw3gQYpZjKsd6ltoij5NMedSx4lbhFYyaqzBa7yZv5Eg6ykSCprGWQzpXmF4lyA
xGyenxEl7Se6+M2gjtGnLpno+1aOGwyQt+Heoe2GDwUM6UEKcJh8b/L1B2rwQ/DGQUefR0/mKJJi
TRVtBT2SCybTiWkLajrABpIUAKdkAKVMn1C6Et7KwVaS7FWg3TA7hKP6GQgiu9Huj0fieEWF1nl/
73RXYK0jse4biYPsEMvmXaXIsFlkZb0M1RbLRAy0S1UDuSstWla9nVKyWjO6YqkZplOEMF/RbmeV
t2cmz7PgGqg7e2nmGlnSur5aIUYmWyUpIaGyvshiafrvlQdTjTWP7nfx9XfOgMxWdQawhj3jiWE6
frTCiioUdHMPFXd6YDZuHDVM/di9W61wUMmhiW+ODVULbhSQYA4DOWBgDV+w+YPQbIb+CFJ9Cn/q
hDzALZuMOisT+9r3QRIDkKt6f2ITNK6laq60CFKqjK1KyEgZBRnRJEdtUoCFZJpURDidmcxi+VaQ
TDBmx8NRgl62qwjmJJPtTAVjSD8o7ePEmB95lTw5tW1KzDx8fVktUp/aYmSjVXQQMrGIVx56mg5/
DAs/gmC6BmV9H7sHpSKtVvpDe+OUvOLsmFKUnYN+mt9fS3d1gEMHN4j6jPJfjaTkxTZsMMtBW7Xd
OT8AzCpvQm2JER0DKIt+7RTrhc47O713dKvvdapWUZ1RlTZ7vHmxQr3iGEDDQzfOe88koMUzqBY9
PYjOmZxSLegSj0NyzlciUczh77rcwMa8XYH716OL4mafLIc8xHcDAcrGY0R82MUWZX1fkcpkkyZg
Ka7VDvXXNwGTA9h+RPDAoj7tepZEtKDNjmH0dtS2u5sz9QiM0pAJQG2DO4/fojEXMcrtFtC9jNHG
3ZI4HWg1z2tvUc1MRgAiPCiAIh18n86lZtkgMtfmf/2LEwX7D7BlRsm97qJIdIbS5u6hZrFUnMKd
f+Mj4OjPSTormubu/3mXI6VhqJvQr7JTEGbHxk8EEuwGrat9Jymh+nhKjcfUaZTmlgmieQgtDtD0
QqMmhjuHlEwwrzyawvPhRJ+KetGMpLvjUsphCrkmrrSClKGnF2eclvU1ebbcwtwvikG4vKkyh/N5
sJrzlVacdkcjVsF+b9r5ePfB9ioRGL8np+XzQgEG/eAr01AUjmYnyrIlh1AL80gPiU0Py2hpbbq6
ptbMMM5SSITFb0TiVo+FMiP8j+Fl9Kj+t+2J7RUjPmJTCC2r4i/LazjAh1t2mCtrX3P8JdsyPNIJ
xn9zDB/xgpMx303M+MORmwuosx2F94bFq14uohU1s01Posyk04XQfNimc4Zrh8mroyBwU5Tftq0z
DTfhqLHHVUeo0Fb3tPg2NnsIYgeigvR0nVUJEXZG4OJEMRyi3MpmSx50mKP+K+B6LAHd3Zru6iNd
7wVJDEKph/jAtYxrjTdeZ3l9ra7mNg4rFa1LvDCV8Aokge9kEIOfLgdc7OtWfQz6ojvm0kMWQLt8
MJh2eDIe711WUnFkvQMfVVBt1NOm6AkciGi2OZv42Ax4h6gwwDiFOrEQKpihsDZudlfFCWmsd1P7
x63Id77/QmK4dwtJL9XJVjBD0e9cZVpWSHI58B4KzgpsF4B2AvwWMI1X7ckgMFZ9R5eku+QlU6gy
K3k4DKHnh1oevxDxabTnLxUJ6094pSe4TValG8tgCeN3714R2gjZUvfOkUK0xqBw3qxycORvjtIv
/k4jeLp2Mil/8zFDIf0tn8NZJiaOZIbnrnTvAwqw+XXLNzqB/FCBPOLeHggaJAGfHlDUIV4wm6mk
nl3Hkj+sslfSNs+zQva8gBX/H5gED5AroRu+byH3vAdbK5ScjsnDqyw1CwUmMnt/CtcayIxiPdyp
tNyO4EFY0qR1COF9MU/YKhAOVn/PyVly19o79o5cCHjAB/jh3Ax/rS6ooVguxIqaQXIeNkoo6WWK
ZsGj1djl1oAakA0ckY6dyPUcutbrBhqXtUWb5JrZWBMPZpU0gVNefpkLeFOgYM+6JlDyhBMXtzl6
lwrrEOJCqKOsM8hc4zYEZbvtVkLji0t1w2Hi4nkXwcwvDwV+hFGfMmh/nujS53vo7MakWT9AQek8
rnEwWAkDyaAlYdwCYKW987ANSrvfU/tQzSq9B6swSIFHUurWNYj/D7jOjpDNRsxhWmA2tXT1bM9n
b9E+tTtICB+K+PuS5nUfYwZ6BKIC3cn9kfHMkPK60VCyyUh6JgiufFa0IBmyQ6Bke6For9ily0zB
jJxd1JQa2gJTg5gEwmq1UvkEfWpIQbycd4LWoKSbqhjSMRtHFzmWQJh/3JcVVF92WCA+T/RD92wJ
ohN5QVjUggG5ix5GWto+dB3bhBWzyXDtXpAhqr/OIa3IAY/gmn815Zyfh+CWm/g1vROACQlshGEK
G9NRGE2WTQsJWhtMA6bbcwtKhMj689cxHptDjAjcbR18lgamsvcz4o+mGTaGj96C+/QtGU2FYR83
5hkdudyygjNBswEDMZg+GGwaGnog1OSkBEFUV9J+GaqvPEsoquEsiji5nnTv/f2SJsupC+wK8d7H
YOJir7gOYJhdt/yxoNdv6ulkSUM7Zuv96sRpsVQfIAr89yARJ5cjiZ+sBnx5KgT2mQ5h8tq6iPm5
pjIG/cCQiMeBdbg2HmSqTSfgJ1wqQnS1Qf9HxBjXFkgKQ3ItvaOOOK9wBH6CAN698/3gvSxZAVRY
UGHnRwU3+fjE8Pwf/dGe4iQeKyUU1ltRaKqHv4pOtupSY3Eq3J5XL5sJJMrJ+x6MMI4lEg0nFmzo
5Ig6t4sj7E9B2pWLRJyvdJAdWy4HeRnj4Sk3H5xkfa1uuQ3XUhwG/bflCxCa9OeEAAE2ziOMrkBS
ugBqR4Ll/A1RCF6n8MlVLnzocUxU4q7JCRP6mK/b6w7vNFm10SfBfb6nEqO+FCALnaUig6ZIFaVN
eif/poiqYUHgoHhRpuISt9CuD28dyCg4dSDYTNbv4Q+th+nelHNJ/fSwvyQIhUA4RjPDFL5MhRP4
D8ChVFbLIui6RydEjtz/n//d0LAhAapUSltsZp+QavO1HIB1IVx5x/c3lqjxfuklnSiXmfspZ4Au
FtvBqFQ1dbKeGoW6QMcEHciJukpJJRo94eV1j2yKbHpAqxh9Nv2pyUyNyNmOsmHtJBQHnZyGdpgv
ajv1SktkHAW3lpeXAhdRw+aqUEBivfCsjuIlxrhnyz6ZMcmvVaTw+1tISCVyemgQJmBaTOYuyZKO
oQ1GKNvrRHog8MK5Q3rxQ9WDePojbKAT9c+iayhlLz468/kAbV89k2/YDpsWo7ZAzL9Eb/x1yGL7
vA2AK7rM7PqAriaKH5xZRqosfR+4nKynj+S4PPlZyo5d0fZBloHINnQPIxGTAYm8/YJoBTg0r83I
59FVH27hdXSUjpsLhVLHBM5or3jWocDpcENOLn4doNo9tfHw2a+xjI9lk5o5UKZDoT2mNwJrYh8Q
g2mtgP4P1Y3IpjWfqo3w0NYZzzhefuSKSaq2EmPZuIQ51eznnMJsEqEF21BOYWbt4wrpEB15osF8
7NPqGyNR3Cto9vz9WoA6k2jUekc9gV7e2va9OnDLnnlQJUA/sK0h9dowg28pkVTfVHQz3JJiivzA
3yPo1jxCz1dKGTzHD+1sBtmM+lmxLYvQ4NDlqV7pGMDxbTuQ065MyVyP0LbLVlj03pfmNGy8ZcdF
Z93SMNz8Xaq1yb988D+4vqH22p7XGJvT6RCdPhJ1rptXlRthB+68rMX1e6lDlgFKdLTWFykfGUxe
Gl/sdPykZahwQY0m6aiA01xFM8G2VJ1KfICvhsDPBhL2CDJUIt155aZD2nGoSQvkfPrGmblTIkE4
wVYXVFbDgzfr/bIQxDB39XrInh/3XoCGFH3WnGLpOM7SHghvtA1VXGn6+O8nVaxw/BsLmxIv8JOK
OjNFxl1Lz887jXmuuFmZYxi0K+Qu+9ScWVSctHaZLKiJGe69dRdM8h0DiHQEefR1+ykrDaUye3YV
UlTOXVjXyHc/xBt8eqEL9i9jNBUbqeP4cKwUpPG5Lzo6Gs7CXl/n9y7A47Ub9uuerpQhctwwdan9
epjHK2MvAo1NlJddbBr+AJB+XqQNf8Q2HxhojGGrctWmmbD2reWq3/vOKTg/aPBOtbYXU3Ux+ctJ
H6SO1rxcU01BPr6+a6tz1RFjC0CwqEhhjlAkqRaVo9wiQpWD4sp5ta3KsBlCeQPeF0eCO941K25W
M8D2nHuRA03BHJlVa8RhpzUSjOVOpha4nxTrf793f17MXdJS9zEpyFlAELouZRHVRB6xi63rHd3X
6KrXZN8HNplL5HQOyDVLCig4oRLoKbzJ2H+wqQjZs1aXH5dn+a0vrdIS/1vxEYOOqQHS6JAfnhl6
ryvW/iHCIznRloVXK7UWcnMWSreb2o4x+U3vxM/pV+QSRY1F8+EBU8sK8kzVm5oykcqmXbLlC+pa
2tLCZgrkPcOOD0Lw5gG/hpmm57p/PgAGasRzceoJ6wfrbOAowjzLWoTVK8dzkF1Ji/k2JiAiDmAD
kQ32ZZxmjoPdY16gEIUOmZ7KSFKgQT+IP29DSIA8nSx/WMWFS8vrRTU/y1RgKdF+JH8R3z1J9u1Q
LefwUEUi47RJVkvwfR3LG7disfKEIjHJ1y5EaCuRvmM/1lbZarmzxlqUvEALzFxCd/LYCHxOzQjy
pMddU8+n7s36hTQIzk3JWNISxZTm+e0dw06xCYP9SnBvTImFA0JVEi4LjFDV87M+MigDzk3gX/EK
9H1juE8OUl1bQN+HEtitbqGmCL/R9HVIg8yISme6quQElbNnCnfk4RBDXnceYr7GOefst8hgTgEO
nEyYmwBL4UrWaFJ2XKCpMeVlVQy1ZXvZYOZuZyOndZ5hqaPbk7pC2WVWIMlrYEv61GbKT0y/aVFg
piK38Fgrb58AkkhKg9YyOxbcmx9bXKmd3idyTfrOJiZOOHX0a5TOuSael499uxuDPVeszvG4AkF3
lkgqG74G7eS1FRsuKGmVZhbReMk6CC1Cl5gJljyJy0Uj2lYgzJI26nuNRxpcShSAwuAoSf5N8ZeS
vInFpVDS5GIrnO4cba1pG2tSNnzj0TPa0QrehKprX8NrmIOwxZ2TLwX7Xqgb7KKVVAvQFDGwiLEf
2Hiwq11ttEg6ruKug5bg3E/sNAAOKxI9lHUGayVb1oTZ8ceT5mPxxWTb+BfcvLAmNEadCf236LYv
LjIzAnw2JbjfOy284uTRlyW1whYZqqCJfTt/U3l5tb/aWc1Ccx3zykFVrFKCpRtmvA8HCiUqwYvi
sPiQIHwjeKSIVD+3IC4cwc48TjnB4lRbgpolELurch8uwoII0wqajt3ysXYsw6r13jeA34ZFEK5S
wNuE42rUVlP01PFNEf5OdF8wUc5w1KbBBg5mBVBNK1AoywrZGsfJzaToq5K9h/42WJGN3xvENFCD
u5MJIk7rR/lQ7YnJHQmbCRtlctSfiuLm6Lxh965XU2jSq0HnVwAQRMSjK1Xt8QuUxyLVPGn0pVxE
MbgyEwuertwVnQ1+vTB8W4KuZ8PV8vKtGMA52ou7700MPNEhbsz/34Wg9LAxFhda+2ps74OV30fv
sV8FkRWqknvRfSSOAF+U/i7ePiEstCDOn3fjKT1LBCPowBy/6d4RzuBZMTBTMcdxbIFMGSDDSlUS
ritHJauMfjDvBqr4WF+PdhGCFet3uTKe7wVOdXfxAOTEvrRZhPcHSgBBwLo7pEUCDbCuFu3XpkBd
g+RK7n9ACsOlUZB1CWfpnDawxeKkoAVCoY7MxrHsMf6Y2SEEIAzSKDYGgtdEpQ3K6iwc6srGjYEb
YeFUyEh6FgX8k/VcI8iKQYZYj6ROjDHc9aNv/19RMPp2ukxNgQRi3WcfM9sudw3KYjcQZS5UScNk
Bitg+gwBR7mzOvAjcxVEjf2VG4A6wN9/fSlzjpUlHHEvl9urY8FrZQVWxkRmstgZuu6TahC/2+1V
Iku7YfG2Ut8VLJR+Y9BYtHFj5iLwCvXNnlbS4Jo7eFIo/gz9LmSrAnrlxPTQV7bWjPaCQcuuUfCq
y9xFjwpc7temEh3VpVkNDTiDYdPosUjxsv4raKwSNqKgmcAFGTX7s006zc63hlon/KIaH0tA6Uo2
McfpUoi0wt1RCo+xM2HL6ad0Ix5UXK6FW40QqrktD60Y8wOKLEinxqpY/sZbUxl8kOlDFT9w5YQf
hwTv53htK7fSX8DbnxcxZ8Oav5CXR3hUnApJJAy9+lL4uxXRXibav2Q43g2aqWRRsqCOwcy7isI3
HgRUB9YzJcsWktuT/Zsq/tQMyoESpQLVniI6B96nbPM3swPkx+t9JBRAyj3m5xeEhmYpEa6OEKCk
PdYPSDZjcA9H9w5BhlndoUbcFYwNkLewvMD7oOLcOM0ba6MKkBLzXkWPS1Ig6dkkxyV0rsNTLyRq
F16AuyZ5qJA2gXZ8CC9MUFQMvEB8LEfjVYsrPbbeVwuFs31ibJhAkaDkrJLPGj0+bhxNypXUYf2K
tMwQusZ0BblS2qM65QjLjiWcXLK7WLlV4UHj7IywXMBjvQyO+JmQBJxtavehAzPP6Frg48oqJJk7
fCx2CHVu50B+4gveTmowTE3ktfTuGgGXom2zJDjJO4yfl54SvN2d+8K5vUSjNYpU4xYHS5mRg5o6
EcRHHM/NUAFKZF/1n+BUah0ek52QV3QRy0im1G8Wzjj2FGF/AB0glerCGfoDMFTIhvdvUDN5C+Vz
rlPKaHDeXQifS8b76R3EQg9uT4VzhLbMtPWjvPwiCvLdI0mxaQTv0gq6ICBirZwPKEnn/Hp3LrZs
V0P8fVWlnO6K/AOdTLQm8Ac17YbfM3yMlk3HzjdevQ+6a3M7SOOc/ljrwAFZV/dtuUh1B+4hwwIn
G7fTijIeReLidvJ+DnlPo1K3n9neY18t9zVjcqe2qXm8RclJts6fFFw3fCiHv6RjJ9ZhHk+aoHJt
EIO7L22eEaOanSvaeJDY2T6w6V1q6wxckzbr+O47daC3jdWSxjKT9GSTxW8CR3rhM+cqEG3H2uVK
GCGbaaLQlcfyELz3GAM0Y4zNMeftjUTtbN6CHP0oilF5I4TWWhCA7XjrfJ5L7KILT0N/MJG49yYv
8J6teOy+nPDIs9GmyMSAmgNROalUJosJPJeH5gJdEHSxD0to4/5qRRpZp6Kn8uEPP9Akm447rVNB
sNbLGqd6UChOO6w4xGVOdBWT7/W1q+mGg7uKFM6QV0FvmEpqWcP8JOuYV08AE+mRLDaf57vS8t7R
RYwVaYJurXFKAq5Bz+HhkQmEn0lNBmpim55pPWYx/bRDYdC5jcqClZJ5fF2WqXH/XARorF3X3kRt
H3arsJHE3AV4fugatOj4GbQPpGEomUxwHf8APbesJpQIW2/qIf2N3du9mu8S2dJmtMClh2B6Fydx
XCMwnjdUYkknnjCco1shBWL8f7VRBv+L5f7wOumkxX6JxFoGdUO+2JOTFv10QxIKVo8ZhSqWBGuF
Z6Y5Raia6GgnF1McdK/cb94JGmWJcriZVAYi3VQQ0b9bawf7SqVVrgmi2FnAZNnwZRrq12V8WUQv
8BXOQhei2dOAIM/CCvyg9kv/Hvc4KRjSyWnjbMGFvAhWspBknnNiaU3BbWZnDljA+e829Bfj31KJ
A3P2m6ko+ZfJkrrYbWv+34w/YLJtLR1qcwfECOXz0sR+MQMRp7BZMsh2RlyprSGnAi27rBWOtlzi
1DLubwk+/2aNhkEUXDcPf0xYgiOek7p5LGoTlrRmjLqf2ckWvrYT2vcKNL9JBI8WDQBNJrAoRZ5z
EN3rszc0d0DLr0NOv1DkM3VPLEbxNmJN7TYhkA4Z+QJpAX0gSlIwIUUMOvAydvvoOzS3UCmaZiuj
gfZIjrDd9P3EU7IIBCUAOQusS8jPwBFU8ny6DDeeKcJ+exytU7tCHHnv0jPIqzyxnQxiVNWpfWlN
+DJtbVVM4Kg9Xtf8+mvWzODNW7OYTtrAWy6elaKjebH/0bNz7IoTYGdXL7cvUJkDRgkwxrTuib5U
Pze6PyzlwXYBkeO6UjiUnXov+2jEkN7N4je0KYqKMs+6QEiin7aMwuU5UubfbZZeSn6O2X8SitHZ
HuFRVz4hST14u0qSRaK2vcYbQvJhGnPujcl2jpT6WAfAcQV9HBJnXeND6okUzONWw9W+qujingEp
fSWJZyC0oCAEPUAPNlMKke6Ie71c1plAusbewsm0wkpmrwQzPYqTU10lZpsewwL1HIsQGunhxjs/
r2R2s4nH5NuVojbrcEC3kE4Bbh9Vr061ZyFs4OnOP/zOSjj+muU3Ppcqj/qcH+v+54aeAYwhMRr0
d+ezqwrKM8s7RS0djUWpg0lA0tny3GheEl6rM+JPJtF2j6bPzkDp33JHQ9LJ3XLnFP34b0dI81vy
NvzafPoMzYb8XQuXcw9rxXnKLiHRZXoKoim6tinynxy9FbCELdBGnKFAtD0TX9d2wmepSQ0zcI77
1yx66YtEDCwzwjDg1gMXGOovuiuA9CNk+jTrsNwxotYyD+eYeG95KcPLQPS4FS32EjQRHmlOxkrd
mVjRGKRd9DMnYNLCxUCz+ONpoXVwgd8Qtqvw5D+v/PkxIvkISf52Bw3MuL7vrK0+P2hRdXc8Kmfa
6KNXV72wN9BT9vcMe9wQNQ4rOPHBBrWOFHrHb3pdFoUTdsZ1NGIxi32/OFAigZHseYkOCar2BZoM
fuZkEotPZaJNS8SWFXcxJzDeAPOTrnj/eOezsVerI7nNhabPVco3XnJri80n4CrJ7pWr5fnfHms1
voLpcYfZTF63Sf7n1LG6fGjpvzNOb5t/cDszff9j1kQYB+KSqJo6DOhFfGYiaHPo5c2SRonm20YG
kIt8+VRIALKuRa8wscdRQxxcUokTe0M6MkL5OrtpdEFJK0qrrFYUz4aYApaiUqOzO9OicPmnHI+U
Jjj0YT3JJewMdWvd8znhbPZJqdZSCyXqcJisTaMS8s7FghtEAbNGSHWWwRz7VmnHBIi3L+dA58AF
msY5MNbRLT/+dLcpi5qIoQxsM2BsjLM4OooFudMRfJ7f1SJGc9Ybn4C3b/EOOEzJ7cD0gYKU1WNc
nWBEq5Qi42EDlzggtZDrZf703wAeMjVC/GiDATyeb0efw09TGlJtd+QskhkAX39x2NrFkI8V/t7X
Go84EvfF6nnY4aQmvVmPlIdsHoNB81gqYHPYwhwA7MKQhwE9fxGcvuZmxnx7As8N1VRXRko0La/v
hK+96uFo8fqufW6hvzyHBLKL04xB7muhRHasUmL6RAPbImZeuyHBH0shjo8tQ51l/dpUqgqudDpg
HVlPnt5o6+sexdIUUUaT1ZyD33M0c1GT2c05SFyRKchjZl/0z8SuaGzey1Ja5lOmPBQ+ep9aJw5k
he0Se55ChgCQWpsQx47ZCML9sGT2FXjygmhIiuoiMaZCBeyYUaN2ts6BctPrSDgh1YpeCE9Iznnk
IJtJyFwrSpTQRhXY/SiaP0UjX/ZnZmXtkaMmuco65us9S2bihw74HF4pv4so0cKixYG4koDHjnFi
qKqIkpebjZmn8T/Oyvty3zohw7o8TQLcDECLMXvWmNhf9ObGxPQHN/mvDHvu8YKamTqRdSypNQGn
GKmCApxoNa84RcV7PBR0YbE+TiIEvImvgSXBjOPLUli8DP45VMy/9TY5QJYDM4i7dQMCqbu4x2ML
7s8pBVa2nLXL+k4Cch10UA2WVc/1yUyppnc7PdZAqwRSy01wbjyv4DL7E87YFrP75ZlgQRh2UdkF
i36EqjrSjMtpiOoI4GKImH7PlHKBE0Lh4PK+a88VVXpsLYS+LdapxdV0x6msUkYsURWoHEW2KEnL
XQeRsjOUHkaEW0qWelztGlmoZLC6pFHH+9tamh9IUPv+7+uuX2i6YXK1jW/tDBkh9Cs80uC67Hu3
YgczvVzcE3rJDwXFMJqCWrlg7IILKt/r6jXHYoq8K+ThMmm9wW2fmSXTtNfwhawKbEJ6azUBMiGr
sqIl9eMB3To0IaSMLKgTWl+XyOttoLJgglT8GlrV2SZ9xhVYzl8ohH5ije7wplDdK8KkBSqCR0Yv
ULgQ3O7dw6QA6Kh/2vSfjbzGuGZkbac55nn+2kiTb3GzDteidygs5l4rp+P2VihLn7y/LS4WuSbp
ipLj36ZyhxU2UC97WpcAalR65yTzjQnUOh43TM5TDfuhvL9bSy7+demaEaEMikWpH08Hw2Hr8C3C
y+hh151z9g4ZvFjdYlQKI2uDc9AfA4OaSbdgQCA/uoWOAu10t9zZAUyIl/G9RdhazwldUvftOZx8
qv9K1jIL+c8BjrBBlaqPfcKgrM7nQNYmp6ELgSkoHF7yPGo7XSmE/NFh9ZjmOKuc1NGMf8wY+Fmw
DUc3cjlNkJeGW3RTeucnah0WymCnZWvuJ8TuWYCPUnudqWrknCtsKpNGvZcSj2yjFGuv1aQWGDK5
dldLqflenybMazqjYLA3IGHRurCt6sFfVI0D4Al6GwwVKhdN17C6FFcFok7vMQf5hc/q2fYgKDuF
D+FECgkeDw+JgtayHmv/hVkNS1k4cM44rGD6im90+tlGjAzR64D2nWKIOgQyvPmtc8aDnHKpdOyn
fCxBgXk0cspLrmYZ/uJOElv3tBWj8iWgtVMqzYBiBWJUyTBF4ThjxVeKJGAkjEJv9ggSMYYJr/Se
HWdzN2U/6RhKBAuHqF0/pckX3KmCOpxOOSLauw1ijDJMHHxxmCc3/8UzVZ2mMwOC6trSxadrJ8tJ
zNdj53Kwtcr3LVUbJ5/cXnrjbwUnCMXmdwyqbcSYjHKSLtdTKYQvoqOadTGoNScELfhBgCVf/usG
s5A8Bdmek/+4mI6osLqjjRpCkhRQjYywTVA7JVFYkpa3NPiUN6Y2gQQEmVHpNHdKZgS70iVNl/c9
MeQxa0VPGqi7OwLjtl1ut0DZ68enzBigRSni9sgKFJkAMRR/SD+S7+wwix6Sy3EsmMrUofedlddl
hDExKw7b3ccWrOmav3pw5jNXfwjjN/AmQMp1Lsm4IREDqcO0fYEd8ZOTFl/BI+aVZ3IdzzbVJWKt
ppTIOE5rJfi7MDSCdOUZefNwMt3EOjHJz11VMttG+vUEuuUXGd66DEpShdDtQ06z93mZPybsfmYE
f2fInoS5hslSOe/V5aF/SxGn/AhCZ0f8v4ui9mxItp7+FIT6EBchINmDzYEvnvskMXlm8qxJBJPL
ImLXojDXJlbGxNDRAzmCJ0yG0yfL3OCmukwMCgf9qigG7vwtbk9bk3nxnSyWD7ayxQ1zM856M9Ve
Oaoh7pPoxNcPTtjY64y0xKQ+bXyp2peCjMT+xJ/zwyAF+1jWm6A2z8J1zOu4rx7+jWjS5fnhGVXA
Bk+EuSkxCo/1cqXV/ozjt1sXliEkGQ2crfH3XBNqLOyrIb+8jjpN4Ep73C9Iy2laJzpNs17t3wla
GBdsSQDyqQ+D4BqUBtLBZ/z/J6x3vG5fmfZcjVC/okdpY9LuXwC3t/PannejHIBwSRBt26OvNgUE
NNDtUsXNsdTHT+cHZXqqGL28Zv0jBong3vyvJnbu2HmxAkKShR1ZL0TMLx81Lv5yDi2FtCcng4Ec
1Qr3a+I1FKUGqQM+umoIqCowhRpxgFi24OPijYtnZwYNCDCos425CQqZzLeq/KuzcD5aAheN8P3w
kS7ShcSN4qct9zzDHnST79GygapfBwk9jNxnFQvbzFlKiG6QG4J3NUrhqjfYrQ0hptagoNTnas6y
HuZv1XNQyhddwMzn6AmbGZ4G3dLxjkqi2v2AGscYOvVyfxiDGI308MkzLfa4Y2tAwH3GlioHdQQr
DLQTAboP8ru5RG1+R872cvnj09HB9kwVD51K16zQy4hYD08ykfp89nxXlHAm+LVXclSu5Ik0gZGg
6L1AYojfOS5VYLdSxloyHlRH9XN4rIZsxeRGWthgncNx9OpA62yP52DUTV8bKvr29L2qD3pRTb8n
wSBQrpruHEbB6xaCEsq4mtL8mVDkxhk7wkRyHl4drFTwnJK8SJf0q7JjwUS4PQDysXVN29diN8P7
ovsrkf40gYbUzOLXlo4nxM1LT1DsteodrOqduTihm1SdQJtuSQUA/23ha+xDw4wGyVR+NvDc4su6
93L23fQm73ACErX0v4fgMqAbHL9+XsMvL68fuur2IotkfU5zc4E717A/Ve2f/jhU0lV8AMU+gHg6
UQUbuqEfw5N1Sx2x9UYkSVTMNgaRGrt9cZo5BlQmAxVVhAM7svMxu7MAYaB+iAoxSD9I1eoiVkUu
tURjtxwmfpQOD1fz/7+ENrqIY8c86w+1D0bLMz/pJbc9lEw65IhYhLTmcsCMHpYMRmhRPNifAslN
w4a7WuFhG8WzdCrp6BnCkyLP2uIWfh2Nj83bAVf5qZqmjekvm+9mmYT3X+ZLeIEBYKxVdfxWWQey
njlkRzMLYmdY+fmEbHMTdzpgI3Yb4bKPgw3drzcg0mw6LvO07xyqH4z1GuZ0g2Uqz5x9SoGKXHXd
QSLP+KaP75KRWkb8peyykOK6mmqc1D8axbD4St9zYua8EcGBbfbjXP8tdsL3YiyaadmhwxIMLnXx
GdFE52BIBv2A/AivsgESdLFT3FxzgOdE0i8nSlwkBuHXFC1MPvVMfyGEZFkXfiEezok/4JFiGtnl
6g4Ad3wHeaPNc0aTxaz7g0DnMH6F8374syVp7Xdgs2k4mz8tehOFPbJCuRq70vic+wzSfBiKkU3q
pkC6tqoJuV4lI9fmEdGeBEFCiNa0SlEjyt2JEeoa6qE4Y+WiA5NcY/2k6MlagwAag4qNOYfmbU2h
RKQ/8kKE3k1k0eTR8WxC32df0rsRMalC4doJaBZc9dMbpuXRtmETQQoYNrj8+mFVYzHo9PVm3V8L
neQL09FnVPPAJat57CajeKOLc1orLzmJaIHEFYriACM9UapMFB5D+y02ZZ1+a5RB6t9SUZlNMVXh
SQfcXFRBWr6pB3NG48sNUNkbwRUTKJistJOirAcVFXtAP8lay3Y/gZiRy15vzsFTzIHIEXhIM+Ab
sc7K18keQwXAJxqs+tFOGl82CsV1fO1xWALEsdLzknqg2ZsT3hrtcXYnQ4XfAtU7+mAO3rOrX/fc
g7sNjzLRDKNUwEt7Efcc9sAeAM4xM+vaBMcipmQ0rQQt1VYIgDL4JXlguUId7DN19EdnMHIfTPyU
R0oTqjb7olUpDUqikuMcAJ0UnzK5yQA4suOJsP07q7QMwRy3J6Es1xaukOC4jK3YMOfFVjC1Q4e0
1QE3LBhjs81SjJt5Ioekz8d4ruqxxOFJRfU87LtOQTuyPlCN605oWjWPHJV4DF59T+MiT57MhKMy
H4CtTRM99Xpf6YtJaQvTwC0zPCa9AiYW7x2DYca3W/rAzVwDHj5opiSG4VYIchDi5fVIzTuVkwA2
RqKI8pJ0qENASarn7V5RJzfPOLKE6jXQ+Sqk5f2p5ZEb1qS5vcWWJ96OTasowwYJFzBQL21xfwnk
hHyaP/9UmMQualwH638kGt2f7bdSkbFXRjOlK8ZJZZUbYsqYFXYX6vKqoQl7Q3eJ7srXqvvwku1x
o0j5uWD80Myb87kZyba3D3x37VjT/7cHVolwYkMShgirQ+f1le962gm9+CU79MB39LUTsKmG3NqV
Ar8Gg15StsPRg27vRiWAStjsfmAo6nzxLaRPN0TcbbxDv1zXb+nA4djzypKwowfppudW+mMf9zB0
BTiK8jSn28g9KYt7qrEHHTRukgDG8bqcEoHHX+G5p0C2SfOMsXJj9ymziORTlLSr62jrU2HjIUY3
tbxeCa2SbzLYBR/rU5HTwnW1R4JAWuJoqNt650japbqNOTU54x2uu3baF/FAqz8J1Oz8VcMXhbbW
kdXy+UglfcENrGA4kG0/GdS7oXukYWsHO0JjNg7BrOd9QLOKWNlLPSp4JCja+q5oU121GqAXToO7
KMKWq92ZPjNJJLATb5xqLlNuAV1UYv988tAOjd4jRXMtr++0Ehhbs2DdIjT9B5AvCJczB/xHkzAU
ecq1h6kzk90wNyZhXHp8Wj+Ih7nBoB/zmrv9lQcU3mU2wtlEGnWsxcbX/96Cjy2PdLs1TdxdGaf8
8Ypz7dnvMRqKAG9vxGMVRMCzLu/wjtOGLnt65UlIcSBS/I+44tNtlGRK84+d1/myL1GWZ6gRdi6Z
OK6MgvxzhOTqyJtVAZbOqHR9B7AbI1yJMtc23LCgoXJKrVdBGsXngnegUTSZMo7lzPuPd6Cx1Z9d
wI/T89fHk4aSnVQlSBUJdZDwsBrRKb2gDV/8eukYGYI6dC0g9fI0SWRoIKGgCX0cR6HvUeHtmM3P
ifEW1nXMyCfbnHy03l6sTPSUy1xIo/v42zSbx/E/9McP7S/cCODgtiwQCt3Uo28tapvpPzy2iwBF
ECEQIM+EeUJ53tPEdPi8oLJjtliDSwdlN2bI+9ifUKi6lBq3pY1Zk5x5jESWSQUZBfm5MrQRggGp
0Ik9RmnDZ3jomhFDZbc+1znJitGhSl1Lf9zCs/kBx0cQ9IRZUG5a8Vjw3shYEWm6oRl5ix7SqZ4U
S157fgIMGWvOBZjG6hucLZja9pNUn072hBLevWPpB8CiT7zxVotxGwkK3cNSfeJpquULfY9OMGc5
FiLcgTSlMXGGcQSUBPUQS3ilKeQMzMgRCap9Z4HJVW1sHRTIq1FAtHDhDNJvEQMM0M65+b0SY2/X
vatryYxyThIIsOfC7Q+vFWnU+WB2AJFmPXU33UwljzlZAPZs4YUveHcz7Wr1lA603CJhbADUHZKx
XF39pzgIweJCMrdqHo6rTVhdQFIU0zZstpikQYJrV1jkR1JWMjpWGatato7jykDbjWKaXpwBWDbY
nbVsEocCh30nV2oxYN0bBgBtGRbcDnvLv87JjBtKCa9CLqd8tfi1HLlfbjXkTdtVYERHQIQrFZHd
jnSHRXc9xA7sa1fQ1TuEZ7Vty5dPVSzcOAUkKXOS03HISXXJJH6+SzHBbmr1chCwstCmHYoQZRrt
umeGojQp1Mhy8Ii1UK+2w682lNjFJfI35geWEHQ8J6ohFayi5BJ9ZMOzunThRM9ZLcOtGeIHjW6M
tXV29lXGooT6/OLP35UPp26cJT2PmhveUGExxpEo8q0NUCqxSHPEZoix5lbs9rR1Z4szXDWLkKYj
7hCPr8KY2aCXs7vJlGwbcoZGASQqzKuDETgbrr7JGam2cmV+7Phjd591X7euIXM6Ro6WHkBQ/Tlh
FvnMfuFB9aWR3m5O6Aet4UoxB7wh05iDSHju5PB0yhIZKXRTPyPAOO0iV2xJz2d4+nFbZWJb9SAw
ALNvpP4C+0NGxSSinQWnuRLEpNYK5B7xRdNU2hm6Z6agS4DeJkHC2TQXZBKMqAbhbyKwA1mm1z8v
QADKKcq3X914Z2qmrbN4LAYciA4+rioxyKcsNs390vndHoHrz9+oj2tWXfKPMHhe1IBA7w8k6VYc
bRFCpv7tWBUEVc2KKz+XXeHNqg2/J3smoDEytViPaSmaM4UssbxkfFlv7vs5OhqCaXOJFQKYswXj
Vdz6d6tj4mPx8kKNoSk1pehUeouzc8wb5LS6BoTvSBFUzbcGu6ByGT6k/YRAuYK6lp/iWTWK/urT
0NldZaJbviOajtiSULjWhR2CsxNOuO/IWZD+HTuiYZ8iOnmGNFtfm6Y3fnPSAKfI2HNFrmw2jYWG
3cZ1PIQPN/EVCFjFC6RBsbzhXKdc1Z0kxLETyvdXa2oHZM1pzm9Z5DI1it81K0hdhnwXtvjr5b3z
7+ptc0Y1breyhSuZJ2HD2o9UhkHs8Ga+VMc3LtFCMXIQCgoasyD5emex9Zpep4KCdlH5S5K1JxLB
60gLpwfCWpGxAv9fj8Xm0jD7ul4izqOw9gjpfYwZ7CXYFzFbS51r+ZmWX2rB1nKLGaxB4A36luGO
3GGsYiLaFeMyyIyoQVmLU8ZJtYed3B7Ec4aaMw231uZMhbcNlWrTJcNHzaSMKMGvy8wErDj/1vGC
MlT22rcWdbu35ZPMwPnWNApsRBSZNYYHg3SnA/zfPSSNcCL5zzF6Hma+MPUQfQsv5uRUckr3anSt
uP7wCPP14u6SxrOt9VkYwARqtjNkqNC7KrYO79NhLjl0Uw6nNE+ZomUAQvrKa88DkV++gX9Vu05B
ya7gaQ2+bgF8ixB01BvRjM7Sfp17nM55YFeE0vj2HIPn++ZfAP9hp56do0NQjK59sEBPAWJg0LZ6
Me0ncW+/s4Fd6NUX0EsGJRgRkPlHnhMt/FXYRkrWAn+wNj+92FuVu4ZhF9SKH/j8fpVziB5kuWjr
fJp4Z1O9KSwwwE9+NzQ33Zr20HW+Iu4JF3NdoAkd8rFiDA+OhzC3JBQi7PUnLpROqabhAETpnSpF
AeRZ+FX3fTxC9V7EYL6mo4SPNvtus1rhlq5I238tX6ki4fwtw1kO6DX49I9E7STfXoUk5DF07X+m
oVz0y+vQIp/yOBLfLRh3VmhRM5XIc4tLoF5KebaSmPBH34ONxYVCcTxSzi3VsUOLfikEpSaQWJ3l
dsF3fWunDpSvLo42dI4XeHBPBrFhE5PzbK7/tHWo5XrYuvYQOUaMEaYgIINYYJXlJI4JpMEhIXRO
gASCztHybGAIU4pyg4G5F3Qdoui1P3Z0Yh0vkzKYElXIzamwCiS2YZAK/qg2qS6pfU2A0bcIMO1h
EQe9A7+tLz08UBrk/0duTP0prTmePaU1zbK5NUAKA33gM400Q9BkDCdnPra/d+VuZbSBcGW8HUBl
B0KXHNYltWALg4hSUSLd5XxwAnaoWP9QbN1c74Wd5dMdhShL8X48GtGqAGU7Io7NRnUy2FTNgf6/
cnPsuFj/ZX659w1g2WRgSg4wzLV4OsCF4MHmh1lv+d9dnwIL4VZt2zt+XBnpRsopU7ux2poykXM2
nV3wHF03eREx0XPFxp9xr+wL35fay5U5QmLnDi38+bduhXEuZPD/N2esjzvWd8TJ+O+CIISd8rTE
Yh/9pCp2ImGyc7wo3C+XJVDOZ1kRKHF+ntMPpit5iwcyClWIXD2ufbuwmET0QX+aolw5y+Zkc177
VaI8diKnlz2JX9ZaKMyW6u5oq6rs1VmXvn4ugMTSiYhvREBsHwiPIeQoAl8DrJxCopNO6xOPhnc0
v732b/85Kp1wmkjw6w7VWk3hS0giRtmHMWCmoD1B/AnFgkC+guPDAyX172u9bWHgPEKkxU/TVTBg
WB9w0DohbJHSdltzGSUKBDSlB+hUHd32AQSXZeU1NXcqcQ6LLMgS1S3ZHVfgVN6e8avuEYukzv0Z
o0wbu17yW6NU9vNAKdqLYj/tTosrIv929hluM03u6PWz7mdO3z0QWVFWx/cix0CQGvl3zWlCCzMP
1uKcqJbalnNStMnH5mFYDIJ5lIhbUqQ1gGwkqzOZ5oiDEuoqqi7nmr2BzKw/HCb56hOZuA7DbDfE
KJOkthEtQl0dWMrBg/+znm3TMDdgLQu3OLZE+WCmT8IYJmaWurx8v0SrPaXrbVJ/V+moSXdcssDP
nE7QtGoFA2C8QHtHv8XqzMHiQ7zfWOBplRz+P/jlK7zlYPLvDp8UTMY2+bESK12vKME7ryrZztm3
8mtDQ3CTrMh1qP3yoeluQ29i9tdlWhk0xxvvw7kLUGKLbMgpOchOiZ14HRv3EWQ8pC1MW/9w8iWJ
xWpMx0AmNO6uaZt+8mg0LFCkobwUtoA1u6lw29CORR/8KjE0xBzFHZVfnKTb1YUwveKxemQ0Fnaw
J21f3SNZtlrX3ZT7H3iUSCK+u+eSVJLIhbeUb7TGozr46JhbtEphZ42VkjdOx6FuAX0hSC+xNQN+
XGquInmuFmuBNIbc/6156Mzcnav0e6fTu0AJofh9SgymudnwUQPOVtmP7hi4lpS0JsZAM7hzpbid
6YZJJAIQjzgZTyUqla2awF2f5dT4NULNBksTmRbOWby6cm8XI0MS3EvhA9gPvem9uYqw+8M6wSJE
F4j1remZA/OaBnmzBe4XGv7l0VQMlsOmwroHscEY0eFFzqNAscTXT0U4lw4zpTzHbQcOKuuOLEXS
JixWk/o5SksfirfZeaxEsM/ayonuq9xy3b7pz7cewAGoHgmlMt22Ld8EOgyHq1VYDpiWH/7A3eej
OUk0XkS2e7NzWVj0jvPf0LlH/OMKfnzn6XabpmRdH/GbwegR7nFrNqC9aKz+UMHofCnfH+Y/E6K4
o/3O3FYi6C7IK/7z9RiR8yQ0HX5BOVU43cdadz7LJlywIM9RuZG44yJWD7M/dQW9zjLj0rZiaCVX
4diH5MEJtVoxrUlAAwFNlsZXbSSsjEwpOv4XIG05p5QQqgUQq/Y6e8CKGGwx81iFUGYwnqty2oY4
Naun+FCofCDbwElGvnnzEvbCE/msi4JdXdk3Nen+hkj1dqP9Pih7xVdM/jQWQT0PZfuxBuNNrb2s
KqcPfHYiT5CrtBTz8MAh8h9Nt0Etw+zpQs7+HRwqaDfxhOfOUOEzLlTy22IZwW1GKu8tpHHlpuZz
ZyK7zul81PxQmIhLR1scw/4LEL89H07VAJG8fgOyqw1HAqzYEAOQDtBs+2J0x8UBfokx6xBKoC/b
szUS90DLLPYz8V5NQs5aLH1hGeDrZQqwNggvWvahDTz+UkBSGucy3V+HWKnCeRAnl8kpbmJuQLHa
xDAwF5lCazhgBP9wMVdLSf5H6jJhdjLdQTGWz8AKfQUlxOkKTs0MdW+bcRXgmPMhh2BWVsw7JSCc
zKn9tWzVAQv+rkSsBc2eH9FU2LriVlHMxzdaohFLwD5XM3k5lGdQ7yEAsGZ2nuahWAXMYxD4ICgu
9+Uh5SyRe6fk8sG2v4Z4r6AY9TxGZRke74Uf7oKM94fMHaVZHJxg0S/f4IjFlsw4mzh6jenmDalA
FX4OXkvMRniQ5vWMT0BVOaEn+KsvakHEfh+cN/VaaQfuJi7dis7Ak3x5Rt+lQdrZEFsAWK34pv2d
cAUxLcQxSgNaNuJr0poW+UoRK3uoIjLclwvu7KJ1kvx5BAizjRcgtDV8vyISnF8LHeWDlwqNCdxK
ueHiDhPBZYxxg9wmUllZiZTqkKPGiqGBNodlt4FaEZBUoCtFpUaK1nkT05hEgSLxtEqZ7W0zaeqc
3OAMBkQ3J7tMR1c494xMjmJA7gTZsmmWEy0bJ3kOwFdxRdIiuQ64v3zkG1ZeQkfYFeEYS+3YjOSC
sSh967UMgi0YWMBMw0crVNC3Q9gmXYJUQbWJC02uxCVOSKXuW08TbDW+ZfFu5eRxoR9l/tLvzz3P
lU+jUF6CgO02eVKnSuUnL1xe8ftQoTa9+sqwsFukY0zdnK6Y92M50ssCF39Ml3JlwAiOVQpgCg9M
aB7MhctRKiZ6bj/MO4v17KWWOjdHFD1LPn9R5v1BSdCMMKYxDIQOxrEZD6UCho6BuJbjLR4/GYYw
D68etT3QvwIQWokTX+esY1Y9WH8fYLBEWfJVOsoYZxJrrtmgURujPhaJYKQ4X7y+Yzgg0wPnOYCU
WoT6ToaaCm0Lbl9yzrhjzML/1n3wTQrIxmh9AWLM0yETu6ql/BicRXmaQAFBkQjNVvqUa99o/xAr
4K6E+DusvtGALJgdlO6RpD2Zd2/o1VK/b1Ak55Mn5pNTb7x2+02KxCfaxVsWAn1rk3l/CrHYWPqP
kmcOv0CdQhheKeg7drNEWNrlEbb6WLjLDy1wxFLhQEwhvjAOjzUutB5RQnmE30erj2rlN0GXVI0T
z+f6yRdE9FF4YaqaFCGCCQ4iOmIKbWUJo6gA71RhflB/xKIjHV9dzLPOGhlFlj+htVy6xKSbxP8F
Pe4OeUQl2LDR/qqzJlv//bbeyPjituhez/+mcBVZIj7xrI1s3gHWM9/u2SiM/xvbUrVbPQIcR861
gGBknOawZb7BpYy/nURk8D30u0EIovRCHCtRvBaLRtzba/M4VuBcyxkr1+RQ5VdF0IENYdtswVh5
oOVaZZ9eVBQsvZCollAPzDxo7kRFR8TJT0DVM9v66k8OCkb99PYQVRoaKe/7noGzlS0ONq7ZF3PX
xoXuzYvm579JpN8jceMqOvWK3ZPncTNiFz3Up041hAr0ByoUf4zcFYK2LHp781863nGD9LkdOyxV
poFs2wI0EHBbBj5m0iQtOsLV2ROSnqsZC9Idts6Kq/5KoJdX8Wank3sXa5syhDoqthp90RVAdZwn
Rnctv/zcJL88k0JXYhB4DGlhA3IuJDjbLl2tPT10bGxAKcdJxU3nog7t5oY8OWOEsOQ6VeUELZ04
wkQlL2PMAiGC/KxB3QqitDmwL6ScBf3gLxhea/LjQumglkucryvxXoVaUcjRvFNd6fvFPUtKzbcB
Qwo+/3Nk8OUz/M+85H3actvNiMUKyO4VRQFQ5VxFpKctiaGFPLtEAIcqY1zNpr1683/PYGD5KuEG
AOUxabueBfXciJf3Rp2AtDEp0IzJh3IrZlqjhVLxSCgWoZcR+aTKOlFVMsQR8DDQXPZ1Ct7ua8xX
SWvjH/LsYS5g/3VeXdEYDQQ8dDE9Km/Bef1EqCoEZzLxe6T7XKbkZhnXE77bf9SqfaeMt4iNCf95
VpFq+29RAYfnRf7peolQddZWqIFjQt65bMrBfzyP5q6wXCV/uELt/NakB2kQj3wwWuxSYT0qpLww
kfYwSNAxGWzMif3PGyrT/ohOM9y/T1NXgHPhIqpAnBDQxN+2sXLXlFO8E20kJUo6OjmxKxbHVzZN
NeVQ9GRd0WNNCv8AsqtRBX49J6hzxNT4t9IHiU7kxyZCtk9oLDM8oFIHbhqZpkyXh1zahbyWMmQY
HdpoT9lb7g3Dbn0Jp5POD3GfvIxXDLEbv1LI97iuAN0MdWIgXrBCXMmvGnd/J0f4ZM7t8itOSt5J
b2jcwFh4XxJcSXAH1jBvtFysp/U0lAsOF8atszW3fGlQTDFjwK8EuinD6NLVENffHWGUJU1mmmli
9XIJdB4/r4gR2/K2jBTa1N/1NWNJ13OJdKW3tJte+9ChxT7UT+53Tp+uAYgNy8FbDnLM6jgFOhUY
CF7Ijz/NnuEo0xaP5CAvOpthO/dsTLAIJ0/fA1BZzkGx6vpRPJTFd2dJEiVD1kxjkLrDgu03Ubhi
lTx8QueFpTMqkH9Py4ooukaBjbrPlpSJJwqSpq2aCtpnKeHdgqjGhwRyeSDw73lYRyhx+oT7/Tmg
QkGmpxfRYESY2MiPDNH3dYMIXPBcq0Xh0bKCG2/uhQXuqz+2y0c4STYGQjcBiDqTpBUx78D1TB8R
9vdskqeIfBc5dG0A+z7zoICKiA93nS2JidE7EN/JW6tD+15f8KXT11b5/us0YPnT9bOq5vqdhioU
9uDNdaf54tPJIRbwZaZm2PvoTVuAehzDrJfEXDE5c4be+MDvXWcgJaOVJJFrHGhmNW6+gJ7+0r04
Rrkw7vBQiJhpIIZLqo/5F079rWFQKpWChz9LGqDFHiLaOcJYy4KmVY0lvByPscYMngvZJZ5o287g
4byw+9Fvxpe0NWFJ6G/3NElBaDrN63O+WNeCJjQM+jaczUZ48JDyUpXE9zlNTEypo6vCQKp0FEdJ
YiG/xnKqO9R1VFj+uKIK/lv2oMgLJCphiijDLHwKWRQ3HxEfMgjwSutfov/8Mp25HPYb2SKjrNYA
0usHiqsBJGQtjXmJnghWaCZMGRft9EpUTrcrtETjOhiOO74U789WUXcwQlWt+e1Diw4lA5qzV6Wq
lH5MlxEniTnEMK0GbEpPtHtooKdm1PPposRi8UDKMuGIJFkOP5p9og9wgUJpv0midtPv25owd80R
birxeI0lUNLSDBIcpDQiXQYK0slO9inDv3TM0gsCweIMLpNlnX8jABmgrrmPObAhP4ljYYz4h9ee
wzjVJrxfHxmo8+gYEXrWlA2NodoaOGpVMZgT1xKCb+Jk1odk4vX0Mt9dvGvqTq/WAwSbzI7xIK7J
LI9WNvE3i0cyFDNyjSZ5Bi6IMO1Bjxv1Eh52J/6I4JdGxgXgDLDOh4R5juod+eD85xSGafx/9rV3
NHHMyKkm0pSB7K2auphrU5Kr+jsnhLM+QDkbLrNSTRA6Mm+33V3esGkDHzfmo+xxZWHxYM9mejRx
0n9TGpidYy1p9I05i4UMRDjuv0rOTggoqBewuEPkwGjK0aoWVWydk5NKgcNZm6sy7psem/sQIlI1
usJgLVjpw3zSSsF0ft7Jyn0h1jKvIusXGMDV7l+zl/kL9//bnmNvmaYqP1j43HnDsFJwiz+fOeaJ
J1WPVbWP1Lyln/oIxylybAIV4LxjXOfB4wAifIfXGPcaGfsFXFKted2QF39dEkPj75TcFMb+/ysc
odhRaX6vdFasppkCW/d2YDVllPSviqDXhzqWQRXN4HVqBccUHjX1qo4NI+xiWm8FQfqNU22CwcdD
lO4k/9eJKxLthbJgNVTwInbYAqbH88xOu+dUgGtCHTGiPmvM7dENpF2Dgt0exCOGWQlOdlUrX4xx
InajGzVI5zrh8Gojvrg6x4sIcHAW1KSfzQVxefbIhod04vaWB/IdFexJN4LdvElv2dzSXSV78Qks
ByF2nEGLA43QzDthsthHileKKNqW/fb1FAXddLlPlUQZLTntcy1/OmqwlvgWGVybJKM+IuqNjP/0
pu33OQJNWAnIzAtHLZSuvYptmKh3uIkC4+DMgBHi11CNFxKJndwVYq1NWnZTdpqegjywHbaKdxxd
SCN7m3wetDEtEJq6cwlU0yDQEVVNoBcbDf2Xplz03ifVLEctjT7LsHnbXifxIF8AvI+kyOzUyDj6
H6P1mOv6FOtdTRrNRcO8+mQ8cu1ZEtOxxeuDathiZrF0iBC/2OLx/tuBLDxh0UpgUyIGZDrw3KIF
rsycVtxacyuEzmSZA+hWw/BQIHPy72Qt44rCKp91IvEA5T3AmPr4KtXmyKqoL/BmkrL61P6IVftx
YjjWbXGBg212jBS1KPGhSlslrp7xw+9fx4SafROUoaBz4gBOYd17Gp7XZKv1uq1tOUIhruv5CswW
z55vLMuq5t3zY3QzzbHsbG8sbwf3mNpE5I+I5aIFyp54pI/DlWLF27nzxVghNRbODLP6+H99WJap
BLTxLoLYFg0jvnft7BpEVCLLqP4rF0ZvKW+tJACQIKWflJLxombj/ukacnRqGCb14Y4TcVBb3qxj
6L08HvZpcasTySQCBKeUaRRK1XjJ3PY4PXHwNHF28r6syVBXDWViYz+ViQ7Z/0Q/IwFqyiYnMjTM
m6XJgks6KZGADyY4O+ODOvIoDfT6yVlPHnXY/ikuWBP7YiDYlodoIpWF0+vqGTGs9/IBSJI3i04A
9eL1I9JcDytFKV+yz1VFfFi/n9ciwF4GSYSijL+9dECOJP1bsRVOS5RCg+ty7Mpw4FND66mMUwXI
aCMzAb/Qfr6zvd6/PWMvpGSpSjYJ0M/9qvQjYrpTpZEno17Y4Z/9xbMRNlqAp8KlzJWabx79N2wu
nbpqhsQVBWLF1clgnW9BrhHfbpbneKAQeIzXGb0LMNQ1UVGMaSi4WOgnhQe7Dx8W/WMkGXAuHShu
NnNeAI1GCyVP8WYRp5AlK+ik/lBDAGa126MY6L4xGzZjxUQtrQ6diggpGwkHC66coEbIKL6d2/rv
14DRkLxJVZezdo/MOxP9Ibg5n7VFWbdUQyX6b0V+P/Wievcn3xJwN+utMSCTiorWAg0u2feERE0I
BBRJBAQ8tSzj3ik/jmJxXKdmGS538LYve+x6Zhc6Rqca8i3SpW4xaPjgm3b+xSxDSOlNLs7lusTf
2BK85BQHtVp50fgKaEvq6ryNz4j6iIGcC5OSRwBUhN9g3tej4QoSp16mSTL8g9S0XIx7ONvE739N
H6zikP7T6/S3v1e1ZN0PftbPK8tvKzmJc6oTCkfuqrmkMnTe1dHprNDqTilEsM/WTCEnSCAnwEbS
tjZDWTRn8E7WX0cgH7UftHyCWh5SDcDMFkwDNa7GNOV8QT3t1M/9aji6i92Ex3OuwOel+Pw5Vqjw
GlKi3KVD1RqyVPmVARCajZjGwFyhe9dmuQw7FT9bK8q2HkzPRHi5fH/n8OUusx8fZqW1CJZJ2078
HRhDB2yHPvz3uK6Hq1OCTXEC+tDevZ1ad7JhazqLbjHGxjUUnzRNxCj1vzg/BnEucHCy/06p7ysF
kgmnptax2jHp57HLX+/dXzjgZsn5aGqbcWFZDmDuf60egEanayT5aI2ErcWd7ElMLTO+0pJlmxE1
WBpa3E2Cbcc+8TWX618/1qIaZufmQIbb8wRzqm6wMpQjnEMDKRwnVqUydD/PIr1E3CZboZP5COaC
PO1wPYV8Job4SvDA6AgzOcHfkzrwKtyAxd6AGt9h8oB377KGczVO+uAxagXXU6YBtjJh78ofo+nQ
KsEljgbyHp8kkKM23nwNNxsbhbNtcChN/r0PthMlpX2SQfPvZx+4Yqdbfj81cZAGGtSfO6y7yjmu
8fp0tTINcbi/HOTL/VthdkXFJzvFLbuRVoVzimsdelictxBYsuTB1VDRb3//AidxiA3JMPX+9Q4H
SVOfsUqWAH/HSk18GYyTiyieCz2A5YwhaJ/AyXYHg73BijjUzExSeLiKbiWIlgIBb5/I2tanQQhE
Kog9nCgxwFp3pmIc7uIXgsDFdFLSdTf08TOr8WIRFJbWuHhO8NYNbTz6glT4l8DaO7mrGVpvf9z8
3bySQuaNGkhD07vL3qRqcxMLokrqkurLK1wLV4d0X/FNoT9AAvtnL9H6EvHVUjZs9gd9aUubYuV5
S3xKO1W8CSJjkqoGOT5ySdC2yVTUHjd78efZVUCiO+benLCnOh426pfwb2/uO1gYRw2P1ny62ItC
flrhYy+6vlEM9qQEBY/PUyPH2WsjpP056OaIRrpCHs1y/oiBVty5Cq/oAx8cO2bLBYpIzSbeVOtl
xichrpsGND3iOjMh3pamF6cyFtaYxUe82JRxh7I1h2atp9DY0CgyX43/5fiUrM12PoouB/XJUllJ
qLWNa+Hs/HpE+3es77g6QdpDysThbZqypcpgH+Kv1bhvlHmMyvrkgVe5Vh7BgSi7zGNafAq8iesR
6cLXbI0OyjKKb5ITj5AxS/VNioRaD8nnDjdK/Aq4YNfOMK/hpyKctBdiNtza7zbI9ZEhlbklpdXA
ndAxhqfsy/SNBDZsiDnXA2vfDi4wXeafchZupT7yz81xL2jbL+Q64Yy/u/3Rzq3s1/Y3/JrUnPhd
s8Iz+VOQqEUVIMWiBJUdIwKmeQPf3pCmxZipz5fMIMq/YIzt83knawduoCca+OgC59qlHi6PGcCC
Bv42sid6R7Mi5oWlByzS42Da5+S0AgnJXeMpak880FGWt9BiEivV+kVac2CVYF6Hpul+8QTKhtPe
qjmWltqO7hi8avA5HR1q91sbq6Tu/mUshJfv4fggnleBlYp5xzzaT1kztzsrf2U4kxKkvquYHpuL
xiESmeGTX9iQAcjsrZhSYztzLBwoGja09qUWsTWHyU4PoWaVHhif3zzAjKcJTJ+5HaULF2CBBuzy
KR65R1XOtlATSAAsXP2a/UKfvTjDHeriK48g2IC8EJeAlFXAY0JFAIOoQlMO4wdBB3JYekOOb6cV
FJEntLJ5o4CMHr6Xzto0h6DD0KA0Tns4Qh8dJFCzQZT4RWuLtrEAplAqT8InTeKsd6Q2nxgKJIFf
pU8ZSut/0U8Ke9HcfzFoTw6rQDG1gzLkAy5WRiDbLCeqqLmk+R4uc/kyEog5DBUzdBM2wmUIhSdQ
Ffg4CgwoZsXkjn3v/bu0SWQ3A22ZiUC3/i89/ZaJE18/Zp9PDNOBh00H4j3OLsaqykB1wHu1qw7T
4RwLSW0ngvEag0K2C9XEa8I/FFsfI5SCJZ2LDBm+woS3OjPseEWZxTM/FTeokbWXQRx1ZLTnCJMH
QzBpHYqclgVPLPx8/RJBaPCIQ51phdv9ynneR/RhyxvS7qM2TBzlYPMZcixnEEuKv1VeXErqFA97
Xnrtbwj3eGpmHkP97Bpys7KFa20SnMW41sKH4pGybT8nb0dGuyx3UPxjo6wkwQstHgSCiM2oJxPs
WRAABDuazdb2RfqBOc2rIylhiY/1sxF2Oduw1kUGlpQaHDxlFVSzWNxPqXk1jsiuYNQIWpQWj8Vw
IOdatsFHQQQ/rxloux0zdSoS6GqiqOssHfugo8nZCdcBT1V/j02VLpiP0laEZ0wx7x9XFl/fjV5p
ybqhgQQx/q5yrAcHd48k9MtNyoEZzd+OYRtJHaXMqON0mFReRWOQPhpjPygD7OmmFkCooP9bYSKn
ZBaf2jmhQljeV3MkvVeJAAR8pJsEpLAT7Ghck7+ED0lNuXT9dTgXCjwI+YB2zQEzmauPIY1SNJec
0BR5wpesA0gwHBopvsyfCEloMkaMDuhpfSJGJ6BW+tOj/BPA6ujcCtgYNVDuN7CG+N9LMgqYPb3J
Nb2z2ELbnONvL1YLtChzFf1P8/MHWL0aHUpDzlcfFlX3aKDk1swmPsp//UaXR2h+Bzm9BlM+SiS/
W76Y8lSE9EVbgS6MMPivQJB3IKxCFGxuQgklIaC/guMYKIbHn6hWPGAF+4W5nh09iGot5g5N8ivw
MARaTBedzZwIxtOD2YC7cI3cFE8wgcEbSyMlJcwbX6v1D0NgA1e6LU15v3LGnvY3us3h8opnIcEy
kMdpg6v7f9f8lQs5iFAvFH3rXqsFRW9MK+uRfo7OPYecOBzqzoW0vTwQUcv2354kf5raDRbysdMl
MLAexMHUCMxLmYlfa3Yq0G9AoC20Uru5duTGuS4YI6MVTubtwpfp4hbsIxxybyTH/+ELwP+XaGSK
/o3DQ3Jt0NwOZaMh80ViuYzQEVsfpDNhW7n2vcTv8fV/PaBhTt0IyeCo7qDiXaNF2spsIEbD40J6
6tj0D5qUlVcgibvlik5A2dvuh7H645zLrJTcOqCfIolGdWoz98QqlSX85QRxClxRO3x1BwY6f8RQ
CnemfDEof0U3Rr6WyIwir9pGqg1YsGloUcy0G1VO8Bn4BGq1DELM9stTi3NpU0ta1r35S0GdfuCN
gs6w4vE2SXoQRoTR/+qIpfA8efiSL27P7Cbpu09te0wum3yUJxdld9DaOXKaUtGZQOvMgoqoFMyZ
yCceL2FQnHC6NZRk2+5JSYnGLA6MOx3NrQAyTT0LXs67huK/UPiCP4pj8rQFwZ+FvUGdHERiA+2E
+rBeIl7zR1cjiwIC6XtUY6XjOINUGcd/d8hjh+oUL9Gw7fdl5fYnAPDHJtBS2LxYEzxPN+p2Ov7U
9XhuyhRMxpNudRve4uVNKVHSGcHS6ZvJECwU4pIy/wLe68WKrCelxaK0wk1RszTDiL1YI9A03fbd
EsxVJZ3K7dRr242Ujg9znfruwpaCZqEsMqv5i//3aZMFNadpKLCyaz4w/K0GieMJdzPyStWkUrDU
PWD1GLZc2XhmXmyjqWiLaIGM2Pre/Wl6UOU5qOsdhtDWt0tmskFzf91waJ3oDn7+bCZNdQszzIfl
HhGSNpLc9TJ6eDc38Yk9H84JgBo9huuju6+FNIYCgkx7XERGYJC3vwd6qpZPcr2a7rC0dH+JmYXU
PVPeoP/AM3wRgVND/cxR5hJpDpLVB4Qi8UxtAUJ6uVgOo4N4XcVY7qpGb0lDIkvWMwNghJsqh3O9
iWlyjazG17QrEy9PQmDEnsGbKS7LQp9O/3xy+pvp9OK4IMEJ+xS6iA5mnzz2NCnJD7Wj2kgzKGg+
KYNlW4qZFn3ONJ7C+gt9CWvJbykaOcYUduYjs6qWQKZS3266l9o2gbXkDmNAAsZNVTkhpSCQ7cva
ohs1m9jxyW5Mmesw20OSCiCXTWNzG97tOmRh5uWG9+idwO8miQvZSuaA6tYMLlEu7Xts7QWGWziP
Feb0vv3+pW9YdBA+L9M/xyRvPpLClSs0GFr0hGu9sBoLgtVyHo578LayortdFt/phAQHrh8sCxS+
kc8zX9+b6eUqhUDmclWfVzERtPFPcK5DGPcNy8f+0YTCbhUHXPbQepHbWbioPdP2h8o1bYbdICmf
RaKUXfYD71Q8uFsACBzuPB6bsiHzFIPJ6nBTVHE3qkpgIp8sdqNqplkZ+x0cp14MpXFWBfVd0RR8
hrcHtlhYwc+qh8hrVR3xHUmUwaGoGDBe6+jnJ+V+MtwDM5WcOZG7IQKjl7oVmlCnYAIu0m6UDtU9
LnHuxjOih8M1fb6U3whyS6W615NmT6ew1E3chjGAj8SKCU6upcjZmvjwKVwFzHpxHesMDr/5fHWD
Zlmu7z+krhZ8j7KbVNhRWV5bMD1liyBOT4ogt2P2T/1DcRKibrQ1DSihRk5I0IQMKenD6Uy4XGYA
KFqsJ1jDSXMYbZUM1fbwN5SYlK+xgg2pKRphWXxoRqKwJ82CB2SsToQ9sewczhT4VTXRqQloLOW+
zdEFsPifhv2/dnRUJvFOcYx31qRlpAwOv6VhE/oZnaZHSSwQHX30mac94EqDxssM5gS1uZK6ZXna
ODYJbUEyT2xRHbPyHYSyWxQTfrsaCaGZuCGnb+aJvtn6w+/GxTdBqg5/BiJ54OIHzcJ2HL4D91Ss
JOoW+JGlhP9VaoUSgU8eTQOAaK2jQ/kLd7eHZrRvw4jySx7gykRTCS38Kaf24UNJskbIg4kR4QYn
6C8ZlkDTx1FtnDKU6gyvyBp2zdorK0MeYta8Eo3FSqrGhNrssvbG+7H57SxTnBaEqckFaEoT6jZa
Ld89VCxZkaII5bA1B08Rn9ChEq9m4a1dRM+8UtswquJNa/jvY39N/6VsWq803QzG9SpQN7AeYQeT
mpuu0CKSxQJFHO3nX4jsAzWkNHWK4Um/JwrkPTO9dbJHkv5TFzuqAtTcS3H7WyjvzJstL8ieANyf
pBp17J6tK9RxadhPufyGoLkolyGtb5Wjf6k6ATie7iv97IDs6sanZeDQ7jrA3paiO1qDQwQvX83L
R1C5jgNf/NZSXAUWWhhOuKrNLQnRqt4hoXlKqy6/Vqz8QafG5T7yfgE+UIZdbY+MA/6Wxxf1knGi
nSIR975Qz1Abuf1u6uV5JLzD9vlN7vsL5/1e031F1n3t53ZuUsIa7/BA8Li22oqeUs9PBuRXQEmw
VGTZwYp7yOXVIbkE/lxRMXs8BxrqE3PSy26f1ns3Gy6MzZAPhsvPIFbv/vpBgBiEshDNHQjBTfj8
xIsYwqfUKFjswTlv9d7zTNJDyXKJ8hWBczigI38MBOnL5NFmO4WevWC9zFZPb7OOQ11ymLSMoLuO
CrC6Am8Y7E3yzXWhEXe7LR9G89sKGpzmEaCrg5KIJQoSsEIiEDOC9q4/4EUWu7xeXFM1Qmd7OEsh
JX+fMcuQZpxPYxB3fCPB0YJOYTMbAguJsvVVKLeNbSfO0nnzkH46haZAstdm8QJQynfmZFtMtt89
s56ICqs7OIoFAesuz6vb1kH3cUnxtA6vGhigop7ehiFi2RcGLTq7lIP/vRRyqUcpVOfpYaSSRM8t
BqmM6BsKaBRS+NdqVLxbH2Xpp/1OA83aUmkix/2xiMDYl0NG/IkwMl2DejmRfZbWkgQSuB1D9IU7
6zZ4GtULswbAF6gvEvcEqTgYLfnj5ZvivIR6aactpeH6WWOwkb34jlHYLxH7r/sCGXgd1epJ4p/f
1vEZK3PvJvHy5a0sGpSjxkcoLx3Sud/WYW+Fx33oy9/e1+UEd6rYvhQeFhpZDhCST61gVNAOgpNB
lqXZXFLEnBoY7ds3Wb+4DgVPjwSHcgW9EbSkts4qM/7qrqo1YhUcv0b9CvFlqL6XZpHiCqYOvjjg
WAPrw/Y7SBEh+socM/7peaHe5yuiFvj30VvCG4XW2mNHM4ypzqF0hATPtShytpo4PBn5qHgbnvat
bI+d//6tWthSw/rX8DKOHvcFq0c+a0DkLrH2Ce0jhQoSa3eYs+zmCf1zOwiGR260tFc3FbAn9nIf
eDzyMnaVkAQBVka+qxcYUsmZxOtclMF0De25XtlnRU93MqCR4XkKRqit+6/DdBYH4HtlNFsmi7XJ
wYnyVbLw+NECnxopsKiGx1p4xpBxvnmHR0c7C6Wk0V0hmP5A27Du18hLA4Bx8z5E144kkGpychhU
qtm4lZ80Q/b+koashmdj/SIP7JMyAxn69qgfcPqjaYqEoEXEjdCuYWjLqyB5OD1atABSZtdPufJW
zzWSirMDNIA/40LfUk7GGWe6qp0m5lUcuySI7dBf3NWTdsyLwZ/4+aQ5gHApVWp0NvFPhbDghCMS
whPuXwBm+nBg8Xr14s7icQP9cJ4gVXoyzW/m/18ZMV1UKaIzMIK15TAcvqM5N09Ynehk6OvZx/Sd
/jC+HWtDDQEHG2rrewYpmyu2p5pK/2AQnhdPufU7rXrhiMwRe4XQaieUNdwzNRB/tiZEV+PMXY8c
BMrypuBPbsy+5c8ibf0Rz0OoKr0/O9BSqAkY4mDQdVUkMWkrDk2H9gUt+tILT3EmJ81ecTlDi3O0
tsLW4jCDPsZdEM3jV17v9OCVf+tOrOoY3iJF3S9QZ3HAb/GnNNin2U7aatgwGyHOl7N6Cvm7fATI
WoI+LqhWB6r85pMgWmR1esqCnaxZsLupBHBxdcBWUk8O2qAVx//LmXqmdktrPF25SaeOdDmkQ7Q/
b+FY442NgdS7+vgpfLfEZFMaA4hmnoSX3QxVGNFaIN/+BeIl33TJiA+go6OPAIz4Kf+uzJJ020wA
PPXYuDEFJwjfPqdpFRMjYHUhE/WvaIJXgGqM2crnJf+s/Sd4BKKJsnn8f5s0Gzy168Yu7k8QhyB3
zXaAa5t6cbom3W1P4bHH6AVvgQxMUhcoRXMy2dNNFwL3dRcA+eZZZ2UAvToSWuuUdBjRRwAW4yN9
92Z2AcmF++scITAgc9Ddw0SGDW9Vmt/yrRaOBcsx+3nJl8MFnupmFWtfX3duNJpk5zPh0N8hQ6fp
lqAv/X/geb8DDzUYIB3+Tqlecz2YoDeSyvfKFISV/PtqK1MKqBlX+r95221a6l8rNJmYw7ZnS48L
OaGj+PSJBIZq5H+jmBCX3yKcXBpbyswSnlednYqyPfS/Lyt/tzz8sFEhJRY/Cj56zQFoFsxbnL6H
zsPi5JqmQwPh9Hs90coxNh0G+aGIN7C6BCAM1LTYYVpvJ8Ww2XdMQtbSoUAvxJRTjaon5x2U7Bcl
JwJeqwUECjC52fLCu3x0/g4GW2H7NGarfo9tRCLFJ14FQWZdML7HqW82VPBUThXS9hVV5rX0OGQh
28Cqxu1hJ3yyE2UnyGcWB+Mxnsq3XjOCaNAnlLhkR9XzZYhI5TLC562XmlG+Vd6w/58VQfUtb258
SVYq3/mJEOJpEICfEPxUN/PcDnEwMnketpVFobdybF7fkh/axFxNStjvHiSzJFJiuhJur2y3YBed
OAfZuUn5toxxvyd/asZrzhORtVHrjWUR5Ltnnn49M4+wyfv++PFYK0btQ4xDIQRc4wpEgEwKyVPv
BK4Wttwu+yYkPL0nboDdF5Q9g5q/6BhNwW69DapCWTTN6dQS94+sQif2NaQXdJdb+qg3i4r7vRhB
PCjdpH1K60pnMsPfSV3CfxpuG76vhuV/x5GjgCz7aEj7zqaWYokfhbtlX7C1EmSaG7aUoVlQXZyA
Amn/D8Se6pdGCqLTAYcixHU7LUtUaWRBEM4HUzBZ7YKLPvk5RDwyWFEM0sW1DyvsJ61N+Bgh9fu3
cBMEV1yG5wWtSOVNkHXcJtk1iVig/MIBP1u+tntFHjTT9UVLkz0zdwObKrVcokr09YUWWcWqg3DF
1n2g3OeOq9CFiFtxRdLwdvawO7YCBNCTTZO+rVc4GAho7aXYlEJDMKAEMDyqc/hDkjEbt2Z3ef10
CfeODapx7CIQvOlW/j/WSk0JMdngolNiBCU+JJsvz6Me4gk4uoakYHGm/Gyvdy2j5Ob1F2VQFlkb
GbdOYlC4eJN4pFwXyHPWe07QfIrhAM6BE69EINMVA+rz2KildjaXVWjxIgXzJDk5QFDHxCL5ONzL
b7pRcZuqCS/loaf3e7cwAkCqcTiAO1TEIopZo6gjdoFE50AwozzCY0Ewo2SVd25ZS/JNY5gKN6Q2
vBJ4n0iUE9VBfP8AwrTAj4BN4tDwLgAS/tsm42xwktd0IZishwDi4mRa19ScX7LRJoRsOOpkrEx/
7G9j82pSzprJbSJLzuq1Uujj7xh1DqZb/+vpqt3oXY6kc+1Shd0fu04GtaOfnViRFCZWVs6XJ6Sy
lcFWHxg7+1hSTeROl+cKR2y3c2NmMB7s0VaXnMuccToekews8kh4YuJAG4W9CjpxIEpLou3RG6OG
MP/S//MJFFfd9B+zBJhrTKa4eYjL/TbKRN02tzdB6Hhj4gZ39QTZTBHvgeaKrat/QgSSnrgS4P5y
ubuHtiNPcIwnfwDrdEQUB3VK8wSvw+EvzJWeCRhMXb/zhOa20STWciS0drH+IcHy9b3sCvGrtoGL
6/7sr4cfIQ/2CeB8fKF+pfFuWDSQaMQWGZc6N9xjNbw61UEoSD1tCsMiYiOPSGqVwz5m2j6LsSf4
/9PZQQscUJU1DLGuZDwayH2SHLcoNE4ml/CFR/VV/10+sWj1i8gq+uZfrKDsClZtv/288V0iDGi9
AnHzxDNwaIw1smIUDXZg6RZl+joLt2VzaIfubVlbzQ2r4XWU6p6iScAIbM7RFH3x/+9GrG25tkki
3sEWOBOuiaSNyeMQMtAzntKQ2qH+aHG4rsQc0Toazrwx8KTsc2AooW4OokU0pEQXR10uTUapWJcE
Rou5MnIq/nynHmgMtwgVisLtZubBU4p8rwk87DBySM+48Jn/f/MV5R4v9vAAC7+ZJp+tpzAMckrt
/+YOPoiKGnnS/eidOGxIefpjSR3aMI0PxxYsrdxv0OMvPf0sC+ymxtGM2B2ADL4BfDMgl1/W3Rcq
KvtE07YcW/L9+UPCY8dNyN3683e42wbMihSMxAy4CUFuwEQ+PXOXmwO7JBp64g6voQPF0fUa/bFd
GVnfEIhjQV3uFeX/TSwSzoL4M0RQ0ac1ahro7g3UqKDBItJHQ4MaZ1b75eF6qAGB8UwDLTaPgqe+
hZgbBrGmB2rim7/bfmjr/CR4ecnqKxboVIUfMGZyMj13PiRKHQ2Ky2IhTx7NsD+OGfLjFfESvVs+
tH8fJMCn0p5R4qKYSMnbsML1qCThrjYO7r9rzDlHAJxR6d/MjtNtxFnn95WtJ9xFXno+QH3DgXYg
xofv18P2TsYr29wp36EYKAKYfGPrGYe/rmBI3Sr03EVkk6rhJbS1NI/8Lkh1Mh81ksMlbT+uIdv9
rwzivAUNjrCO99gjYcRCSyo72W02FeV4YJDxU24F9/On/jTGBi3sPsYPdBLVjym8aRnjyQ/VGGT0
j69cavsBXXRJlzr10wdov+CNen7fC8CYD6WIiO1Y2bbNoYDB59mhBuVftF6xtNZAilRW2eo1fI/d
smSZlN+Ofexy5UE/snH4wzT0GXKA5pWLuqpcT9hkbNw4DxiigS7GeLwCOjF7a6ek/KGKLQXJdKsu
K5yjWSc+WZuQBlnC9I+TARsZsiUZDX+5L1WyJ+0helSI4aKYUpwu9Kxv2YhSmAIO4sTt5OMhi9P4
95hXTOe45urfHXdu4qKuyqo0l1cFOApAXfyrvDPbNlbkt8piH+hxT7GhuPAAGK2gEmw/5xBc3Y5e
8DjYDS9y72FsWm/owRjkGoXl3jg3BXWdmnhBuvBKd1Oqk4z9PvSaWNChugIOUkAv+hf9/o0oTauT
05VNMnnU7yJfnuyLmIEhmk3qPmuh6SGmREqGDCuirCxnmDX4dmMPL+NHmQtNS9+JdyGz/rq0Tktb
eOPcR0/h8BeQ28WZjd2+Rr9QOKCQo6zAl2opFJVhj+1TC+RNJ+1ByOY4CIuP3HHHCX6FuS7+Lv9R
93zWGnqiwe6VnNAJMdADspsM0EfhsREG+7sfMytogzbtJ1YNEYsJ2YLtxCpH5MPEE/FRsA7U4v4K
xWlBNM4VgCnkN034qq8Abfr3OEE/1I6YWMeOvhtC0lkyP990zvjpIgJrL6joy703W/QMO/uZKSxU
nIiNjt8D7J5qevuJVO1SLi0XGCs7hXZk+Ah4adZj4ykWoIGYS0XOu4vAO+64Z5+8AWYPlRmV5Ylq
TYt39XXcefAZwOLfnsvkUReqj061qAPr0RzDo3tNpPxl2wSwvRObieZRmpTqxyL+TOx9ASZqf3Ho
YABjV/bNGg9KUQftV4udgc7dRl0aykGNrcYNFWfGcGtAuZqlYGxZ0aAt7L4R/HkUNKbCWWTjWCZ9
IDfyJkhJZNInrjGBa6MxdR6z0H6pkgvuLKrCa9dvd6fyFIn8pM7Y3sXKdJeLo95EpORiQUk7u4gY
+lSmQEZgfKjrtE3ZRl6twrhXWCeQ5pmgGxkgAVRWw3JRuxbWyoOByPgmoToGduJlg8v1vJKzu3fq
PZIjO0WqFlFXUKIlSGvOFI3Dm0oHIEWMIs6kNXdejF8ez5aGDY3mkk9V3IG4krtsOXT2VdhrGoB8
tMXYW2HxxBlemupIze0l0hbPvdmLey2T+lTWkXvL+33qfYdcY66Pl5N7YATjGGySXdvFAAtx4sHr
KEcwpye6nTQUIgSEqIhQwQIMTQ/z95ns5GByHbP6/ZL5CSQLIOvX9FvJFN3yoqiG4ZFGFMgKfdDl
8rXBlff33M/d+j4ytoWh/kH6zSTtgOb+IR92BCxwokv7xapdR9GTDjMqvPzfj30c+aiBpqH3G0yX
8SclBgonPpWb0Bfjo0tAh59/2qBGrh/hijXRMKKVnNEnN1f6tT3XnltQ5sZYS3hOaZdCFMxIxyLn
Czss6xTaZedk3nLe32uqGGivk4Ym0xMddkMGxh+oqlRsCF5uegF40dx8Pa9r+ZTZ+olL3fYG05hZ
doiMnBrcF9wSXn2ufJXtKmP7D2njw2OCkthiVbg5whErRP+VpjvCBeYt3cUTjYGl4f0pgSyAMXn1
XHmkibHJ38oo4WbtFMTgU33pBlV/X8UArmpvYPwU1pYVFKNtAObmgNFS7R47IZgehT8qDxBVhDnZ
xwetnGtB8w+mJcykoJUN13SqYmZyWAZ1CNYFG/S39yn44E+Vg7ZCn0vSB4zfbAFm7OTG3HO98bLr
ev8Vj8PM9qdV6xf4vC/lA/oI5udNSDugnEl/pSxseTNvQkoNbC7Z1ZmdSQjbR5EkfGxk5bCNAsKT
zksKSuRiuFG6t8yvXrMpKrym3QTT7YUATthemFO9gOO/h+9WAb34oOXzgrMJKDqbbo2zRARGC7fM
zXQ0MRWxJl/JE8fMy0kOS6sYW0iRbjPavLWHUVFJkaUqDASO6dxZ/HojjPAWZ48z2B83B5VKNXAn
eGOeAgDSYAWkRfu6FluM21ZeTVBz3ldzWeqxrzpgAj4mLYtFC87dCxriVsh36HYPbG29S7KAW2Me
zXVSvjYSCht6ZJYi4H/SFl+u4cosBI2Kfkd9zLwJ9jFxnvdsGFUa2S3apROiIwUvblZGNUmtEh9m
9BGkaWaxmE5oKNSMHYhcKGRyCK7zwDu9gUpRrRvw7YbeZd/jbS77IlscRc/4QfY71t55Ktr3BQt1
ujXZRu1q8EN2txX7UrUdh/IFWc2tkxpUDtQdlTrHm3M+gpvgthRiyHx05t5QeSv5vrNW9b8qI9KC
BCmaidBGtpJmVB0+xtRLEl2XGuClEHNmOEGCZ/mlsjGl0jG5XoN5Sim2YagE4DS1kpuShmGMLqkV
1NzNttHxOE8JJkG9qytN7yi7QBwyEJ2ippIyRCk7ZDVsgbhb4smk9uuQqq7lA3Fz9rH5vmSIK9Fp
ZpOn62d+EAxqEyWVUvMwdRnjI3PCauF1tWqx0JbbEYeIawNiwauBEL+z58jL7r6s1wsQ1zqI6N7b
E/kd/F6GMXtamcexgJJRwfLc5CcjSEHe2+w1EfyA4BAdtBiHWbnqmeXCeq9x5iirYr2GE4KSrdJW
jbZSrZtqJi/PAceEpBVcve21AFAZcFbn7Ap5wSHf36eJjUui0QTEEgFFg/xiBg9Lq8UWEir8OD+t
NxrELMBFDw92TIFVtY27zUp90YvQF27eMAbimyq1PJTZbGBdiKUTr9pcDKjk0V4UdCcadMjttikw
OxKHnQ5jypCVyibDOBPeEfSw3hq5/sX3j4GJQqff/1Bz7hY2SIOCQro4uyguTiQs1z1hIdiMCMuk
yWc5C5MUo8jLdqJYANZyINreGX8NQXfTYxRyoMpB4Gavcet3pi2f6uwmKLr8KRxe4xC6UwfWRH7d
/ACXJenNvDQTuOIBtcQI/ajdQnGJvEwsaG7BpOBb12/8kcuhHobdupGpuE3uLvDswW3GlW8NYarQ
tqSIhOQ2KvZBbptv52kIrf94iSvoaCyKVXHv3AzbFbOdwAwyLfaXhiF35rH5YCj0oC+ycU9dLnhB
OuGQVjVKJj7GgsQaQeRvcLV3i/x4BCGIbFM9fjOJKN5brbQ69/ZWtqO/WpUVXFCGfN4mxEtUMnwB
TSl/pgX2JxBEhDD9qzm5lMHbM9zHoMfQ79xTHPX7uxgBliwrJ7ii3JDg7XmuNTnd17kZ3boDdhZh
g57EStxoUmYiQtSZWmsh7vNXOZenabehAmCvF8pyAVKi9+TTBIt/WPJo62+y9haePIYWmr6hK27W
l9zmAK1zhHmeGFE9dh7Y28/xbesReAsFrJGXB3m8z5y+ryEMJqCEA5WQI/UOsqRbwa4/iH9o02Fs
D7W2heqemBZ3KKNGfnw9yfzAWqMEkry9wgYnFmzH5I8Q5SwzQxXmeAaqGD+KlNOxUvjuMGzbVc0X
4zmUBzeJ+Eda/uCKu4Yt4dLwFsn65mow074lnX9ca+cwVyKnaiGfurneyv1MGCjqppYLG5p9csQD
P0hcwdHJdK0iY6wV6xZKNTlgoShbIkBGztfBrEuNPXNvJvjOZ3sLJxIsYtq5l1K1Qsmq16NzGIIn
lqMwAC5Qb1dptzP6dW0xa1oMb7nNohffh765Q9IkCJsJbnjQ2uU8cKxydSFMfTS9HVOO1BhhpErL
GfyUASo82486dTqeE45gV6x+noKXRurv8aEwxbQIhIJZd9LtwpQvg5VFp+leN6n777oeKLKNfdas
N7PLBNwGEfettBdRg56Q/YoVwBPkkHsEQZ7awJi+jnuQJuwqKEKt3L8bBI/KvZEO0w0V76EQEE0W
nJEJZwaN2fwPW9wu2GMSQ1MbPwRr1I+kxon3kri0tf8B6R45JffiFrzD9Yg081PNhxB/lHjwVmPN
lVSrcbONb2wayya4VEKpjhtaIGieiGOpfmnRB1S0yUo77iCH0tO/0QWin/SHRozN+Gh2eHTZuGKS
zTwYFRidwVd17FsUMupW4Q1Axk3pjcthiS423hMxaDaWuPAgZ1MtNy4cpeAxkiF3jX40S/Vu2Mwl
nOzj5scIVaj/6jmlpV0j2yjJggz4N/m8HuPclrh1NaGaXKLfzUfCEOxmkkK5VT/EFr5L3ufRCzYk
WSrGtghwrwPl2aFCvjbaj379zWKkJyI57RMXjlI6rQyYPVFpOAm9Y5Zf3rXiScXSmlA7PMRFUhaM
WCU1R2UNYa8XOOv1tsf0185+fkXG38jvnN7ohPG2e53VbUCKBygH+oEI5SBRC9J4DaWrYvpzosNo
kVOKr0x1rmbWb0iCXaup5WebGuPSlsz1aocWh8xHODHarE57V9oy0XWDUCUTyaeZnEA7yI3Ffz6J
wqCdH321Fol03+CMbENsKjQVFwbLY6wzc3weTQDpfCfvHouNeBliflA+vSIn2xyy2IekKBk/+L/f
s4Q3it1xNxdpaR9qlBAoSp2mzWGawHF9M9o0RSgg2Ii0GUZ18vHy79YUSTVh/hkabvyIJa2inPuP
5sqGrK633QbFN1v7Mhzmfy9PbveTs2etAywngDjNOjiBkGg9tjzDi2GGoonjkdSNwuQqsuOqtJvH
Mw3r/jE3TclAR/gItGH93MrbInJwbqnHClSQpVD7J4DsIk7Yb+Ka5+bHhWP76hZ3/QEhulQHRmaP
l4Th3aywX6axGuhEAHul+TnmL4EGOedH5Jk0Q5uFSXzF2Ms9xOSZSl+eivOwdH/URUtbSdWsrRKy
iwy2jnNw+eDNhdXjmYj46PwOSFS/pZopdWD8P8gU/u5TogDeRUd0BQsghs/xnFsUsk4hqj1Hoo42
tat/+UMzzxkWNPqisagY5nqRxoIXfr4cgfmVw9tO9IYE0Sc4cVCU/fg1beRkGnV0yF5FWCRFMvGS
REtYcwBfqf5Drc/e/BiCKnbJI4O6ZfMagMxVqhYl0k+TwvBzfPnCVas9Ah8s2FZyA0ihOGp1vIgT
Hh90SZS94GufE/BDfFhiWzzlIOMH3buCI47qvtGqFU1AMJFpJC0N0/WIpocsi8w3apS6GQGiyZLh
oP0fbmUoopWmb1Yz4s9G61sHsMMjiq0DVODCDjwNAQB0ycSkfc7F2vjbrEYb9T36qkZOzmYEafs8
u1leP0cKqyk9++pSrUPHeEFQPcnIx1/Ga9Vm/1ZNUDVH4EGu7J5iOeEDmmHpbKAgGhlPB4UwVXzP
JL3Q3pFtk5KjCn1wFdxZYhfgboz40p6X7mmYVcA/CJWVQeCva7bl0+jJdPjq77Q9JdIJ5zrqy84k
n360HzlVakY7LX95D+ARKxZ20kqqVzCMHRK4Wf2kxONTB0Obq2D+kjKHD2vsmc504s9vCpDwSkdr
8lQ1bITcMSBdJaRSXVIxjLPJ4oHvzPnjLXbATiPFfv5+ubNWr2Krb3FRsd3+8hX0hqEFWJQVmOAB
RCgNCQEj14bdvaqrwM7ANxqiC0ZA8ocqAxrhXQZTiQ2IYu1r9Dp6IhUMdSOfHZoe4YdU89gh1YCj
dmnLpHb6w1m6X36h2djkoWJYS1TepgviVWe3FMOArsnl+plnF/QOPL/LDbs1iXstF8bTphsCqbXp
CndgB2M9b1KqcgffJst+VHPJOZVkbk309TdWbM9lkHlXfROJqTGRfhcRiu1AIgVkWWKgLy7JRByY
v87FbAK/7FMKpwFdvL8mqBxvyxY/JFR2vhYfhU0J34BEvRoctMRqAKTJmMp3GnAbch51qEfN8+9f
RVFEh9+DNtpOreXrw+FkhcqNPkLpFMn+SXdbE9xDq3guKZU0xwb6nsWRgDe1RrEZo9b8TK0+2fzs
MKpDr59XVjJtQ6Q5U4nBRDR2Y3XOMFszOHlngyjXaujUOiF5f5IkROTC3QtCdjmgrUqnDykv7Ltq
MhzvDsb2w37NymjKLLMSYqjS6B2yZKCEZPxeYQRmPcrflG8GqSrtJsELqesY4NSeF4B4YnBvivxR
2dky8KB6GlEthfhnfD31rAHGW1nqs3sNqEuqy5R2sRgEMLbZpURP2QYYFENskr5DoMdln4r9KHZx
8yR/CqYCQCVhR41B0w7mKkT3d7Fjm11Q/HLN1hldJV6jJljCebyyeTYz6wNThyNTKYzsU/jGypUn
ASsc9GB9/8G2Bm7VLcygJG1IsJgJ+yf/SxkMesiUOIjNYV2ZPqqkIsdR07d5ub2++La+g3zc/241
hSsj9a4Rg8DwBi0Vl6jt32HIf5Wpd1kDdB2qLzIAOQziU3X5Ql/clCTvZtzvTXy3rpLdbgq4t39q
RqcDhHU9ZiAnxj+BKb8o5v3uQWqolLBLDxypJCBvU0sIqpixzV08WTOXEnBADBqDqAzbvFMyQgOZ
Z1Sv6dQk6cr0F5QNSEaF37MP2q7ATo1t2JPO4AgNIoP+/grSGoAuYeYgbQMnANAr6BN+idUblqpF
wfqi3wMs0lrdna1JR1oNFG7qHiSgA7+XwvV3YGp8cFLafVabypJtDB4d9ldHNBNoomD3KR/bRVwW
vOfDlzoWMHFj4pTdSIEPZBwHDjKMIkQWRW3mu0LLlYIHBi3fuCdAhMrAab97ZUSs3n33g/5HR9g4
AqEhilUP4nON7KR+r0zegAHdOEiaRi8AhNt8coymEKk04Saj6NOxzbz++UvUmrtw7LfJPWMj667Z
KFbzyyoJ23GyTYY5+GDyk9+2LvJKPyPfo7H47mdE2ElpDyD4HgR6So1lnXcFlvpDkk043/J96cgD
5hi9aFQMexnIa0gfYG8tETBybeX6CcPwClmYlac7STgXdEhhDM6t9tlOr4To79MLIoJ+4pdMlDrv
a0uItnhKUnLRmNHYhvR1VmLg3SZiKCcdohFIRNmMsEMmzC3T0sd6BgLGbqBeQXf61P7x5r5GpJUL
+Rt7pvDKa0JBHFR1vZyuZ2vh9k0dv28UJXn94zMAVT38x5xeKFc/UqU+cXOjySN+gW4AP811gi7P
CLVsx7G2TdRH0geuarXJMR5/BnA/LHlQ766OdfLDb0RWsVtL1opQgrin7NmGgnRpvTD93jDkuLe5
WUVzmoCbqfZwN/96Yw9MYZ1SzQCuZd87fLkp9SkbRJB0XO39R0Nq/GjsQzQrqS1n4do8I+KxC2gg
p99C1ONaa4RspmpH9pNEzJdhcPun9HQTvtGJqGM1hW18xefEm4vuhn7xcidBHSIwq3YHWZ7c0C3t
JLkW13Kfb9bbrfX/gUVoeMQa4O66sPBw1+jrTZ/TxFvP8yx8UCnEYlZcC450IBLqXk6IUOqbHLxD
Hry9962vj+uUNJG9xMlT06W51iwtvVqAmcWODAG7N8fSlKOLAhW90RbAZTIE4qhUvIW28VwL0fT2
EOPWgZwwTYf37NQEvRyDPb67VCtrANRifbrpJEeWiFH1zkIgB71uVs2D2tWSIkGWm81iST4J5jjz
aMvqYlwmAwGSAEGade4/yY09yh5s6ZfdtoMUZRpRmCGFVae640FPIKF/ibsVz1S/fXksr25G42Hs
D6ckBMWtDkRvylaWtgeTyqcTMprmTTGXmf96u5y90PkzMyicUvEkI9ZIpU7Q9IEuolvA8it4qJ0G
4WA2SvAWShY5L3cGRpbt1W+KjfxQHghC2opGv8hf0C5+0w+uaSrzo8pZ2um03qr2eAwepkmTxyPr
hxqKKGJLMfV5PqU0Auv3UX0Dru7jpHG2EuSbGC3yQ1NZhJp5TN2dfp9B0n+OctFx/t+PmEZprYg7
rjGhEAmN1ntsrQ6AvHdMdfDdSorR2pPGu0WoWi/R126KybD3dtsN0Ro1utDuPgxN4JcPU/F754TA
bQOD8fZx/yv+xj8lDArY8LJL9PE+CaCqIF7ZIFaewqadPNa++nZvlDeIvSTOCkEHdtXurdMuj0oC
j09xNdJDErPMIWShpK1rZyQjMlf1oG71bmJL7oe2KsU6TY5EqKU6YWyAaFSQ7Mw041hO8eCIPpQp
xfPc14fmchNkPJrcWKjgm/Beis3p9O6k4kptlUpTCjapFEt1BYs81mOBrh3744p45LnZAhi3dOZs
gDvSQRsV0VLPBfC33QIQwrggU/YD1e7oaUNdQAbjAVJSHMv2jY7SNSl8B5BQ5HJvn6HPyXrS7Lel
ZuVlSSkV4imF0xfLTaAXc3evDK1L2hKuGFC4IUxXMyIBMFs4BFj3zTXF3HgjwspISya+763ebLa8
lE1ytnwsUfzcGkTh8G0BnWI7PdPK9xKHjVZXT8XFlvGYaJmlAZvjZkT7Ybu3wzE0F0gkDCc7kis3
r/WR4kooPzAm4fzKn1MVasZqWYq+2U/nSNwmJbqdtiVe4lQdXBfqTPsqAnerFOzqQKGw4KQI22Ny
YXMJXpdilq5PicIKqMN5ykmc8P05H9EDQEhnIR2JGSSxuT5ibxTBjljrZAWYIRYK294LsJyynIKi
J1X4qB0X1IN7WEktf06BufV/IvyagXb742VzOZCzBmwU8768l2jVyBb6jL+OK5oNSIRVZ4Rl1mtn
AbGWPNfvBY5hZSr/sGtbbJWnzoJif7+ypTJRH2vLSsJbLtl/WDeSU5c3M2MEYuXpsj8XIRFI+LdZ
xcWMgY5ihz3JG3ovgHCn4Czg31FAMoO3lLveZXCXOWzuJr/lneElzCBLH7MtqGgqCkkTxtPZt/yr
/BlqjGspk8WfuUQMrcmaG1mzZPK2gXFeLvwa6iRIcqnKuFvDcbbGHMpOtTNan6F40HUtNjpR2PE1
YwHoNgA3EGWBhgXSsmzaFlGXczrTQvl3qnk4L/hclECcos89oRwNAVGUdWgF4PnR0SigicejK6uA
mJRZyIHXBSQTniQ7QejCzBn5oCVJiixtJJNk7+2mhjFJ8zEmRAYkgR/No3JoKU7JegDTYpmb3n8j
gpuL0s62jY3c7dfG+Ro2GigPCiLhSfHfv7V08VQ8QHU2vTT4FiUFk57VO1lEaeojiSi8+qnhBWTV
+xaNRUsZwkAo2q0HHss11Vvdxc5C0IX+lH4d18r+MipFsM9sbo30NG9H0hgHf/BvHekt/YGOpG+m
28OukItpBvu3b6VOfprZIC+i7W7p7SQ8/G8a1FgOH4oWQKXzUlV4u5OHe6vcxmf6knS1IqHhFau+
xdQgJYbomuP2HenyshpqIyqawqIznpTtNAycb/FdS0UO9pZdz2Q3dojYLMqWZDNCxlEY+UdOpnA9
HifF5JxtHExVliD3+GXWcRA0t0RH2HjLgJS0dis7WSogaJWvOjMxs5VghzRuXrFXI4ruokzDbUDe
2JMvvD473bkAzkPxAU3sqhP1YJwXY57G6PWdBGeanSDhlWmf/F3XzYnZzVVBaFqcqMmLxszo0BN1
wRlie2Yi1BHMEAdRAYx+nyySkhYoSleE3hrv/MNKGVskVukuc0lneq20BvHh1awlo9ZlV5hNxxEt
YOnHFD4Nm2ae2jF2moA/oy+wOUMam/dgU2lKcdH0t6PuPq4Ca0lZXnBN9rHjPD6Zw10m0bWdPovC
JE0Amli2LHvikmZjAnWqpxUk344Ge/fJIUdoJ8gSx+gxHfblVYMsSLtPXwPNgzBz442k2umsuPUv
41Dnxine33P3vgbAiglZ028L2lFj1u1mdt9+KbPngtWFYf+rJc9y4dmQvqhF+CSoClwAV9YRU7Fk
D9oH2gPYat0Pmn2J0QrcFvmsZr2KjFT/H28uboe51g4DLLHX7x2ug7FRnJuabYkRxsB0X/EX/AB0
eRoD9XjaULC1/uOgl3SJk7PFW3eY89oO2ulE/KL/xQ5prWOSzsBbmdUKwfkk6rQkLK37bTAMhFyp
nZrc7tHNli/WLjgLBd/hDEPwpdCikz6TpQ8onwbRwTW1tf09JHli265WAZe3yATx6oEDAIepiour
Fxnl7borI5gJR8T9S4a0nUqAOh4q5u3H/Rkt1o8o2CZiNHFhQKTBB9Eb8qnnMK6519V8Erf/bRm/
E7fCuu19AaNCUurAN5JwV2Fuig83X633kJFIT/sMgIA8lpZxGPsTANCCrbOSvgf5EFX2eJuXYSil
zDDKJsHs/j1ug/vRI++Af70FcDyC/VSTC4vZJj+7bgwLThFjnICYZZcq8Z9+giPIIMD+KiJy4MMW
+NCTANqWwDlDAUmC4/+F3O7U3Ah7D03ivgG881er5/FTZaCCwWetjCyg5gNTQFIiSt/WtWArvuWt
N7G3ibeE0GBEIXQa9rxxY7ch8dF1hPR8jx1WjBqNmGmYPBTq6UjI57OKUA2b/05d7HPryVrJoyU8
N7a87wPfHb6LwYaydq4q6xEM/yShLXQoLlnyHrI/Uu0f2L73+TyYaa0/dTV6T0hGzoq7bt2rxqeW
cS4ULYTzCpf3WsP0Tbl+Zfmsf1U0LPgsh8RYH47oCLP7wq2mGTWCxgLpWa58YeJkx09GF1QNtBkz
lq7EUG9zMqYyaANULaiBhmyyhuQ3o4O7bSAukvAV3Q/ZsZPQSli/hy2MtOlMty+xRVmAbAoEEWaH
9KS76mR4FMuQJtYPXsexw4TdKf2mwZuTgf/uhdrwkecpOuMFQJEJa8SC3aw6Hk1cnxeCLVCzBtgN
h1WkUu1CTDr/fyE1upfeGZfRzv5/FWG/UakGHR1JVmF1nF1kRWoupMlCVyR0ComQsygit8vegDZX
Rt5fFY7xq7rsP8PQe4eFc5GBaYncdCnYta0VkkqbLXWWIjnTtk6nVVD5SygSW5Eut6bwoHZDs2Q1
Qya988JlMavaz0V1z/ty6KMVbl6T8ChYGYKNYT9wmA4V4xHHK+oKbhf0gF3ZR95tjYDtIRWSlo4p
plRE9tZ81wfdw/f7bU4sBzYoNb1xgPUgBbD4ToY3st12keb0kv5GVL9Kuil8wMj3TIH9KcOKFLQV
mTAxdB2ic4NIZYrVYHLW+97pr+C1+03tHzVOg9dqlgJXAYNaKPpSvrRxTrKnbO56/aT1IguURrY5
5oCBm9a7Vn7KcPWm3Wbz9qkmLydbKqjteykb47kO1cPmdDJdlO+JQLRUBiAvwnyAi0Q4P9DrV/P1
ZelyFIF/Q8VyqbouQQ8mk3+VsanqEDqGN+QBLxfyi3BoEV4R92nbM9sTl6WkrQd8wR8f55R7B1nx
7tmvBfOiLM2/k+QCjPNwPz6y7k0ToOG1J4gHvETVrU/ZF+AsXGsBGWdozRvoDEWHnCXgvWWn2lGR
D3Xasxti1mYVyFKKw7Yj6RDTDw85Gb2VWZNitxvS+IDZ1juKtqro0YbwDMbDJkMRCBLvu1btLg65
srLafJFFp5rdFNyoeK4Q57IHUw7N+3UC+6L8Syk3//yknsyNcmVbPs+N+XtN2aa2GP8zJdK6F+UB
UtvjsE6mK80OdOG7G8TBhrp8k4gUx5NXYHczo0ree1N7s1Joef/x1zSo8aMShYxwSrgdHN6C1N7x
HTXrAZfafVBCUQfNj8V/y1wOGXdnL/aDbwhLOmr/PCGB0rCltWgUwO9AqyA1v4RysCqoH8pIvdPr
dwlygfKllgzgjhxrD0ksf1C5r2N+/QrFRgZ4J/EsLkXLnOxhYqLsjMneqFe0QsEKqlTvOLAWTC79
U6KfC1iVvR5kBK6onjXrvYtEUUof/yjZs/ZheyfKpgSAp/8zpkW9X2a2TcnjjlVsRkZhC8rJKETw
3u+famvhPS7FRrxVkacQznfQRgN5pVtkuALLF6JAwBobLRmZJguk+Q4cjC520i97xqqSojEiDHZ8
WjLgrwqVrOmYdPelTo381GkiKEaha99AdRqcf/6G4Fclyp8e50PIhfs8j3PawEslfIwKImxx9P21
V0H1TvtDSkEcGRlIGeEVEWLSCW5EhdWrsOiCuoX4KvlbmK0wMF4+2kLyKgoSc/FoccGWFwFXi/BG
MVhJySsfquzmjqS925vqx3rajPd8OxN6JOKnsPjJ0N9NgNMo+ol+bAZ1ACAzvwHYHyfKTsMktN9E
GE4afwRB6wvwWIw4gbcoJyQrqr6zKQw51YeklJmSn9L+yEaTZv3WcIKK2d+itY2CI8ROmic4TTel
RMAgW7nxbZmvVCglv9BC/SBQdXfuOHljok6YyEmYEwmW40bL2LSCEL+a/9FeBAQlvEXAlDuhhKqh
5MSc1lymcZKb7H8Xp+/bj+/nisEtWA01ns33NZBWXRF0V4Cv5qVGR08LkZfWpknbafdmAbMf2M3q
nqO4s9fbeTOJXoGEoGnEcCOML0HAy/TtRyZk7q7vjWDe3TouJmMoDKL68zybeWwSlKTsmDBghOjD
efhzwpNnPvEzZbmrBV0Mr8FHDlWIV6VtynhK40BXc2jyb4JM86fmYEZPI3sDAtI1gQ9BQYsJJ8PW
G22zlXnD11ZDIKdJZzGZI8lt57vWx2ERaP3GglqFGUkYkdOF+ay7OoOD/m1ELFKzi/5/KQwlIzC8
mOLK/lGtYNL63XgRtp/LqtZG/lAseBo7b6Xk2yU32z3NImp4VxhDbpSVS2oXHIUa3Ct9wY4xvJAJ
9M5J10jAJg4d1WSUmoyiwxHqJSS1C7pMOWEEGeFHRUMwrIMr3ZbxQyujIhgD1rpUkFAyOu1fhnMJ
Kfcm3OM79ZTHOFRgYZHdRk4gUtms0MLkTzGdyNyn/m+hnZSxHQwbMbsOoBHsWkFGguyUU+zkOdlB
DYHnwMvugjb1NKIXFKqFwk30MeEAdLZHpf4j9ztTbRrD3TnaiadusvoeEj3+SQRKVuEyQHuO4TaQ
QrplDW/MTpD5OtfCJl0OSNu9tuqMNNPKjYL7i0sWo0q/gJKW4kF/dMX68J9J2MVCp4EtEhpMchqk
GE8eO5CFplTArIfzskkoZjjOjP2sTjiTUjf2kI0qbPctwgQ8YURvaFZ6XPtEKqzPpL1ZyKK/MFHC
r0dxj2orRH9sS1zb/gHlSmApWAPiffuqunYOCAg3R4uhkyKmiV7N/9YESzf7yv7D8qB6UYgzCh2A
97MM0b6CCOKIJH4x5mGVccEMhfzaEu3yPrWUUWl9lAjj3tohHftDTegm62ci/t4YI7Ul4BaANhcp
N0jMtw7C1tf60n7NtC6/3MdqPf/iSVMAE2Isj3nvoUAY8EaS2vPapnjcImTq1D+j65URpOQuA2yS
cnoFvNYS6k2CE2va49WR3b44gvtuVXIvpAnMZlN8kKV38B8PsFULM2diWN6mHLLPLF82O3gcDMa8
AN8+P/5qI2Vp+qIfPvVHBC2PRYUQy/jfpSIpbMY48/UiuaDUBjZbc+Yd+UehVeft3ti6P42LWk4K
FOkhBCsUzWvsJn3P8a598R7xASPhTDmIMGGUY8LqJst7hCt97Nk6PWdzhnx9eMP71OtAJSCGLOzo
PlPlHJejjQBJ7A32DardsoEEEsxym40kdVy6jCubM2jSapWkqbjIwf/4UyrPaT2iTR3KMrXQ10w/
Df6ft88KUj2SXVe3B3Pk760jQEktrdHQjkOoBuappSW1yUxc763Zbyz77dSTl40fwBij/S3znMgk
+uJEomxp1PFK4cmFkedeO9FjF6WNiqXf6CUTgLdIEUEFDE0ND4b5farFtpcYicclOnc0paWBtvg5
kTVXbEhrEekIqALzTBxR/yzmhH5Rqip/MEZIYKEAh2jD541u58Y3fZXN/dEKi3cSeL1FT4G2bp9q
X+jTVUIjLbWjf8ZekIV0eNSNIg3GA75UyIyZEU3anqLoHcT6v3NtVrUsDgd89EDYo71cxTVgmpkk
prWvTlGlSZgJuaaxBM4uZ9CyJ/PQJmguHhI1E4omDoCG7HRYdvE/3xlDVOY4o9dnKjPpFcvq48AV
jfAqhuaQNpLRj/EwwB+sM2i1be4C0G8G64O3V+HEY5NAwHd67lxdOS3Y8SlqIh5vpbsYx+ye29Iv
8kz0h8qSMM97XVzEiCkY2uUJY8W+6wayN95lHPy0/MTzkiyOdoGChxzDG3kLrrPwPQmh1o++jSj2
YupM/jY8sbFz7LAxhThyqA4KK1XK9zf6XwuoTr2ovTSPqQg7eHJQ5RVxiGiuZ22l3zGoiM3vMc3r
gnUe0VPD/pqmKYQmDpdFucb6p6yGPQ3W1lUmvXQk5FBBr6B7GAYA6zqQAgDrFFUjq6B3Bux3YEVL
Ag6pSDau1puLMR360sAI2p5d+uhImwNExX9OwQt9Ft2oty7J5IB1gynukye/+MYL6KpkpXX7DbJX
UsiNjRZp454+AG6wKMqJCTXuQ4mL4iqw4ZFAOVa3Wqqe2sM3IMSAdaIUOyjQdWcmRNMLvD6j2rx7
3jHKCFyK4CmlmjS1tSaSYGoXjGoXbWSCovvDFlvBBpJbJXSH8zSm8s2dnrefsDuDn6lkbNN2oFQi
euVN6qtl8Cxsqrebc/ICWMueDFltP9lHEAFkPHs6TgXl86y7nUctVRZ8RbPpCUXygzqn3MKa5y53
kg8JfDqfXGZcwxpdTWmnCqN5x9VjLik0qpdkH638qv1V/GkWeUega3LHXZU5WZ6g5SNm9uOqPb5j
15f+XaewKPZFYPouang4g+eaPDrTmpadPbIy1QVAALcRufkF7A1Lt7UAcufbQRiCCwnLy8YvpS0y
qY87dM84X3VqHRnhLkLtiUrfNrgiBbrYQilKVyUH53ZS36i8xVA95xe1T5tRSPjtPkdby6ZkGFYj
wSgnJLUnkamonEtCa+OrJPgx+DnWwN2vVdBvXq1PUCw2XkNfNHGYGVboDFjSvAo/ziueUHCz/MVg
CY09Iih5hdR3jbtLFjV3A/6wWcp2SGMbSqKJSPcJXngVE2VzQTv0HACUqetc/oocVCQzDrnwNMfI
ijpnqJtdeOyfvjMkkHutHdYNN5J4W3dOgzFP/ks7pdGEQFW9cndrAhY4WWoYnM3TGkl2mxAHj1Tj
5K0AF2+uRQaK3i4faqCeIZNbolouB+oGvKIVmqZ1kZxgAJA7n8mkJNPkpvJO0TBd1R/4n7gZNP8k
zUr5isgs5gsUuga+GySncyo73tFx5QMfWIJKtjG7j+ATxIEbcxgmNz3jI4OIE/wThWqVgOUKXfUy
ak8ZDqAfrF1qXW5FABfk9Sk3l69y/qgY465Mpk+nQPsTpiV3ieW/Y+3BiI9x3snKLd5ttDttl/xb
U180huRVc+54WjaBX1vyceOrDtx9nrqt6+37d8MmTDYjqKn5qrgqqhjRcFpE2gD3D3MVsZW6RMO7
qupYHPcmVuomz9sqXiZiXRXdXgiOrGnGB8vjnNvLrG01kFJpABahHRM2JHg8QqaUQqw5sszAMngs
IP7qudr1TbblKCKggHh4pZBB7kkvZ2aQR5VBYXRd4BHxnZR1iF9GxF4+/7xiQIPPpYMEs9NgaDTF
o/czkC3eJ/XtrG3dwE8mY8nqTLuGjVYWO+jNKfO9Ba34ItjljjRfOga4Fv+xBKFWa2MAtefCq6Gh
khZCeYkkxn1o9sQR6jJ9odeIXgmCMv0xj6lKyr16b1hKVgOXKlcTIXCpWILB+r/5HJ2m0Z8uFxES
ChTRMUYDhPec1qmONfEZ+2A9QwePwzRVcjzUY5emjl070dPYYJutEECQ4Z3PvvPO8r5TFfK0Kfmj
c9KrVVi7M4XNzz0Q8WjKBLdfF4Te6Xd05mhvPi7YWi+sxmsrmsLJE0xLp4NmtDfuMRP3mK5+kJyE
tSy0CX/Kyh5fVor4blZsf3z39+Ml4rKfNFxpkyaCtGpRiGiO+sLpIEPELCOmCiWNXrWMxTfBxTSt
uYTGpB4GH7usVxFsAj6uJZZWx5zIBjq35Z3NFW/W0yQ1wBxm8pRIcW5U5wciQk2R410gw3SYJGF6
eqGwPcsLi+hvK0tuKgdKmqI1gvy1YlIv6qt5vXYC1WlR0KZEKC/Gtp/tNrYBzn3zQbCrtxG6NxBO
jcxWPCShpXThlgukgfIBaRMHMY5eKsPiTREYkcHftSnTxn3T8XMdWYS9XVBjldVy2yH2gVRzWuKB
BFMUiBDvai5FBjosXRkcQLYe4CIuxm84exLbrCdTLhk0JnMGopjgoHjcae0QY55fhkZ+RMlDhbCT
ivUuUAZ8G4mEIuCsYX42eFJBE+ZioPDLUiJQoQ3X8xrXb7XdZY3OAQRwdBzpub74A+Klr4xpXYUp
NSQOPLR5vlDI44p2q4aqzN2RY+t9XsumQZTjb6xlW+oiHgiY4+KcEMfYwBLmLh1+zmVRmBHF8+la
+/+PoMFmYBInsD7159L+T9ScphaZijEeVH9hkCudAQ2nJ/XjR0RE4zzl+3IAmX3gmffeUhkRPwsV
TEER1rkI1qfZMV6tQMSdIOts8046Ji3xTHfk1arEoWTgN/2nVI+QKq3i1AgCuHU6aV79AtYQ3U0B
vyQfknxUGFQMCn65gZZekfrSDOMzEidKJ2iWE7HQDVxTneEEecrDzUgRAC1wJEJtq6TluVh9cWzD
niQN5BUBgg+nh2b6LuSSfS9YBCzsI15WvFTZ5P8MHPgrY3KaYO8g9Ekusd2063giq23CZfy8OHBu
7n4q88+qIuyex1PfjkEgGxvNY92UP9GfhYwFUA04I6dHCEM9RSG1Xy6yDsXB5woBwfqzTKQthqfW
gC8//B/JRKZxeQQoR8H2HIK9F8ulwFokdBAH9e02S6saDKK5gzoplwpucytvaGMKMQirJPcNUZdK
xVHi7wTCtxkNwVIb1BMWKZ6sPsQ7+TB/jl9Q0dnVwZv6O6w3I5TH+CXhTJl+asuz4IxCE8IDMyAn
XJLK32m+jkKSCPkhmsV3bJyJ9j8jNAw5OyvPqkPliHvue76cHKGmaCCFMZUQb8J4ubX3Su8dQ1Gz
LmVoT3M4s7s79DPCN65J1N2XV5rzzy5z/tjfOYeJcaxXyocMxOqcStrlnxls2WZODPj1kGI5XJaC
QaTjTykNFo0j9y98vnSvQ8ibUHeiUbriDzYqD3d53lufpmEEzEWwbHw+u8NSAUBzzPQHTkffYfTT
TLV1512UJMovLxae4ihs/ro+F7ZwWPBJTsk0GbYAdmnWPotIFVzvrOg32+FJknrtjbI6oFabnHSP
yJoKkPd6Z69R+8Es1jwP4GMyOkv2Oevgtkyfr2Exa9XV1tRKNFwoHGsGBDh5NffGXM9hB/KQzboP
G5HcSfHQAAxQvE5kIY9fXqR+xrss/1HvU4fOD9elml9OiSouKiN03U8NHNQJcQxgC3TRXm8HLRZF
gqjPFZ62j+vGGohN9IYMWsv2wbHKKvrx5qmbytVWeaW4bleJ4tIH+XW9Rwhv4kv/tuSpNG9e3WNU
mn8RzDkre9f0eD+QhW7e9gbgIKrCuwNvyN+uN+OB9q4Ie7R5eOTmRYJfTWjTIDLnKVOsU4VPe6Xj
sfquvPppQ2NfcEEudPNUv+HNEyXPPKYGoZPnA1KLPe4VYln67P9xFRmawZd15kf6eLsmi2g7kVmu
JqTrFfBewWl9Afl2yWY76smiyr1T1iXKF0kCH14wmWIbI8pwHnO3z/5vZZIdj0dVrzqaW/hmi4yp
IckMIr7RIN0sBsyX/euTbdSSXd6nrK8AvK6m1vNOSFz4fkygp2bXCgmGLgX52fhMZK2aCFYEQWy8
GGj2ofzd0qeSaTRk5VVn7bKDsBiSA1csWtdG93WJVOkoNqD1ohqY/ipIYIkXG0zwf6eMLUYzuEop
jt/ZI9pXXgQo0iJgVbH9f6mCNH0PltBsCDJXSxYRoHJoVHvcXdcGmEmp50ETpepEeJ8UrESVd/Ts
zACeo9ScZNxWx9pOpCvYPV7GYDRpHHgI0AHJuELzzu3FUKhHoF4ROdIPUB1eY01jurvh3kLmrLfB
nPbhHrpKsmEpef+refQz3bvKn5pGo8Z3pdcaYXOAwfDjmoCdcruOGlgeccEuT0ik+YhqAMcXflK6
/0P29PMvekQo6RCK6n7Pr2qrau2meiPdWwB5V07CpIwZXsgjCOYl0NQwNnkOAeLRaTsnnip/k3TU
fEQaFKfGOkS2YNQG0RrwJodmaYnXHGHrPd0lEttz0iiRhSrhMp817jh/EokgiGtlTaiN7W8pwqIv
dZFXjeJdOOIr8oA12me3gH3bKzDlcTcEMOdhuhjcQw5BTG9PA1unKkroiY7EPaLj6umii+YZY3ed
ZQ0295RjVypURDlceclepf3hQcFIjqTR48XMKt14p0PjznuB6F8nyX2oS3Rj2lAy5xxqkVSBEqEV
ryCGy47GtSk28YNya9MUkgbHvB/+A7r9+WySokBjr1nbbZqstMOWiXgqcCLPwZAjgrV4vYDGSyu7
APg6czENV0qlo8mUAp+tqYaLckatbxDgRQMr+hl0eGr4EPYViZWV0XJz0RNJQs6XXQL75u2TThFh
e30jHzqChu9GAH1W+NPA9tZAAB1Y4bNp/pz7eA9mMXy/1Bfw2ALLSGUM5oyoq/armoUm3em6Arw0
+NR0TzEXCNmuDHT6J/4yJJhauRmxAiD+ZPOe1S1fJEvq/BE+I/6r7XTBJ1PQyDlit3kWlp7f08aR
5nhat8iIAKf0anfHWiMOODeQlEx7mAgnCvOJibiIurqxMmEu2Lxtq4pWbernkmtLl2R6w06dPcYV
45AwhRopysxBZ6xAomCnZQtN7xy6pN3rqMdfOpwZsOO1PnF8wiCu94c+hnEUZQVnSHa7XpGQbvQD
lBDVzf2z6gWoMhTEVxdDu2MTkHqk69VvdnE9LubApUvblvFUPYRnZwFFfHdjTlRBKVAqdTO5GV0u
L5L3yc8fI4MV6uYjHKkLJa67MDJ89oP790roWXAQO3odQVUXczJNOEwuo934lXiAXW32zNAksv3Q
qTweLsJsMI1ygrUvECK3Iz42Dwt1Ilq+o1hhk1LQL91IWCXrhTsCQn4trPtC2NygFvf4eNwrEcME
LD5FjG9X2KVLTRJ/tgpsy9sIB7ZYKIqys07IAEvl7eSmI1OY8+zsblm2z3xKvuFbUA9A8/cDgkSn
qKqESyOA/2o9y9SRTAhk8zTosOMTSKod7cXUnXuZ4AkWtWdU4IzDDsvWYLs/RbFjjlF32CU+zOAb
vYcA8Se1YnMeaueCqGFi6O2V9A7/SDIT2FmRudrcjUFKx5Ib/wWSKb0tzTlfEmnsZ/PiG0oGZuWB
7tm0Dn63aUBvSIZfIjSsfR9YFG4jtbdX2R9OXrpE2zIyJIw94+xLw9mkE12GIjjWZZZBgxdLG4Rk
lpwk7tyZDD04+lZhSKJtSDKObgUZkgB6qisEK82fa2CvutCaLW7izn+A41aDcylbHxBKfWCDNQsx
AfsjQhioGgUI1AYUyGOGxPEwvfUCQTvW0rkzlOV570HNVh4kSOHvg5uoGfAOvPTmh1pzU8FzUP0y
7gWN7sN4SfkPGXoFKdBn711wtjXfD2TXjrW1Dyp6Tw6cj9VsslsyDzTdddQaLiptStr2N4cU6tm7
qs8GFV4++Qtythrcxx/qrll9PHOV7O/8PS0LnemGHSmb2fhSVbKIKXeMejnfKtyzjL8+Dd6vEY2W
b09QFVXZ5JPUWX1dRM20jZnX4miMLgXcMsk+ODcKX/OoeGdX47233IwHQRu4+7XaGdieCrCt25i8
ObCaSXk7UTiaA+0ZWnQiPIcOiyvOpHKVUF7tJsSad5RyhMxjSWp0qGT3rnNN26jtt0bzE1GjGjyR
pS+gn6nN83e5pWMYlgf/3HdUyX4CNyq9yAworSqli0ax7NCbNtM0oH30KUVHTp6XPneVbFj1l7Kj
wmfJCaOOA5zKNeKbaELNIBCFnAWOHzEjhSfQbN368CqVvucXWs59VQonesh+TYldgVZqZ8PG0fN4
vdkJMhcAGeaPZMgFV5lJ7gBsZOqIVF9XFsJznUDTlxpodl2a36BC9+qoNWtrZpHuzM+PaWqA41s8
JsNqgIUp8u/ChATes1uqqTh+557jBk5kpihpi65zUi/kktw6ACE+HXzbTLxfOuc5H+iXARCmPQfs
PcJHsDFmvZpO8/zEHpcnzBgRY93yDxslCw2nrnxfQf8RMsS4ZgL17UV6JeIP+K3NTRn3lATuwIoy
rUL+BNU01CUg9SWPYRDnv0wtP5wzLzGxtunwV3r1A57gyDeImkTPY/WzZ5xJrjP/3x125mYaol4A
lWvFm2PZUilRRP5SK+dYgMudDaeEVjH5rsfjRhnqJZ5YOBngihtjC8Vaov9DnmBAxZo/7/80rF4Y
VZlmgYk2hgAi9RpzPqcvqUc8wE/sz+hq0mf78IfJqgwd+rK111tgE7Ts1qBZorP+yD5COxm6Hf59
83J1E0htrssmwXLEwXoKBMMmVeIZ2W8ibuNEUabb7mK72CyT9rIPI+DviTNDGJqRQM0shozTT6ow
OEpTIGc3QLyjzsQo8hcJBiSHKuy7JB2x6MKxncoCr3OD4CFY805KCV8O9BW3pnqZi77FkeNZyJqJ
Wy707jmYL7AsuXPpTMb7EmxEv9wX7kRG9WkJqGqI7uyAFrxrz86e/U7rhjgNM3YhA6BRRe+Rk/fG
jekwWcU2BMwYZXXdFJWZe9e+6Uxg6ksnjCqESQ0RdbGLYFtkBBcLge2K4Pa4WYGjz6reF1bizTfa
Kespp+9jAwk5DHyVSw0pX759dx8BkOFc1ZRvUqKNjb30WkzmgTk7CLquOWdHsnvS0Csn3P457Rfo
qcCwa3xFlc8++9LpMjhLohvRiXIkUSvOWJDOvszN3hXdF7TFKVQY/jgSiOM6RMlhrIPXz8ewJl8K
16zNLcpNFIPuaL/RIvtwjPWv8OWg1BZFCp9+xkVGAM1bmshU2XTG145n+kRuqdtpmkckCk+/R5Pq
ODg21cSzRqauCIRZIV8unoSMwB7WG9qf9ij33hwCy2bRNpJ8IVB7C+w32tzcpXzQdV7zEoNMSE8o
kElRtP7a0LuNx8t8genJU1YvQb30z8f3zml70Hjlbw6aAAMSizLpNv5ca9E7QQj+fLI8IKNk0HlN
cpnfYvauR+FqRNu+DS5rTCD4zN5bDJSBWFHY2l3uZXzpraYjs8LzrxyPaRWr2+Zkb6CLvPe6/1ZO
YhhIHoh+YxmR99dd4sY4mh+qlO8bCV8P5vQicmerb7hefntYHUn9vqGEuEN1TBp2P+UrqqPmLIlq
1Z1D4NSNZ3/BgC9LFFWd6bP2pngIO6/eLEEwMUsJNQvyICL1TJCVZKhicG34fdYfTWnCfK39Z49n
CtYAzXAFpO8uTX+lRjlQgTn9xA34UID7iioAI5fMFgaaWmxDBwN+6QYLlIcCxUbnNR6EQqihhzah
DtevujISFmUNki+bGlJbucwZAslcizo+xc1bTSl1k4agn3mLnQmuHNUaXupAU8QXm53w5CE2QqIR
e/wPRcUcS1rw4CoaYS+R+GpATXL/aY5wHggWIYO0iRgRnf+kGU9YGD3pn0/v6jCTiW4ZlKS3Zi+W
8WunJ2pKLjEOd7/OJcQOWmXExHRta2xVYu9DAcDQfQat3z7cyZN3DF+PtWZXGR9MQTth7L+h56Hu
QIZpqIInufxRyWgdfq7evdiEVtzKbPmrD8uhAz4Igzinpw8Z+TKZmUJUzH9F49yqL7nx80Lx5hFM
SdglKe0Ad+nlsigSq2+jxRiz1jPPpaCb8gB82AY7IznvSTtIQC6eMv3Qu0ex9EUnyLcRT1Pvfg/e
OYjwGPhPmhDsWkPoPQ5l44S1AxI5bOC3YqwvFBwK3cDJGrzTnO9VOTRByrFRh1WL8NOwjjgn9P+6
GR68DeXpMhEWxBqXlsgTMeZUvgjJPWC1zC0tDAXVbls+qTGCS7oxsZNkrc/T2Wq037cmmU6Nu6hD
2tzd59UoWEotllHtNB8lkmcYYgeQY9AbC9kAYYBEq1X482PQiUrauXNdOdk/doNACTcZdpOzdnSC
KhmH1KMpkUWn2FXX358ytFmackVizp3yrITALHlxYcw7kpjxWigRp5olWRHS5PWz2JOn7NHEoii0
X1InoRCXO2DEEh0Yt4pwGQ+O0wxqssSAsVE20+Xi+IPRDFdVODc1dZrZDqLiieibuQdk3TjXONHx
rLxd0hqcSiHHQb/xQMVrZBmMKOJOp+SiaUus+AM4ZZAQfjobB0FtSs7Fvq0Xh5ZH/9zg8riMxtDc
8GkUVhFV6THztCDUkNNafQGDiTIInRLbWv7mhbv5ztcOL/Xd60xsW0m0meNLpyy4GRpTw1yanVp3
lF6+sjChRb2Y9VrJUF+h/oCG6JUJUzGURYARnGVjAD1E8hGvJSCnj2a8DJQ8R0g8HVcRlpaJp6XK
kNrIvJtBd/J1Kj7nTc13Y/jBY9vcEORiNJzo8bwn9gGgJCoMab8vuTzh2vt3LCIavtTOxMZQ1Mr6
u76djdbhNGz5EB8icvxyMgLTiJli5svF0CKH2zGe+eZCLy8zmDHBKL+DiCNx41ch0I8bWYX4tRUx
4YWpNcnaAaBiWEeLptmZ8yVSD5qmAJ4aKzriM6DaU7qWh8KFG23F8y0NEBYWGv0+6+5eovM9oTew
orqDoyzsVS4r4wXCT/CW52Kr3Qou26RMAsJ2/nwSuHGU3j05cHjG7UEETvOE+aJVdQEYhDwBpg4E
iOyoeSpFv0tj56LvyLLAAq0/FuWtG42uNr8Qtt0cf7QjU4QHsyU6kF7GCOeeZMolDwkXzQ9w0gsm
WGC3qfUMu3N2aCBW1iQB7cc4T1HotMpzR5BND6dAPEyjhMUtQaTp4j9eiWlyhf46UKJW6fPKyzIQ
RAFzZKLA0qEkedhMIRVQh1sIFy7omvSpPymFRxuiXcCBgGReyczyofjTSSxWWtT2erCKJJ/TKvZ/
SaQXeOn8Lys1pniAYzGGowGYFJve1HpU6ddzt1JPxn3GwFkaeEDoYhBa+Z4agh+NWSxi0iw43MS2
NbevqcVTsgBAyEUbuX6H9sF+HTxyCTQH75R0lUuW7fTvILzKG2xF1ZQyHkkLH55jRWtMV6QfZlzR
7qodl0hSxcO7D1YH5ejMUtNLtSNMzhe34Y/q1zBc9WdS8a5Mqwr+z9KlWULbwIVOo6M4sv0uijab
U8etKyb9mJr45rTbknIraFjsA2V/2AAkBdcCkIys7r5a80ex+vItC4lNRr3VmE3S9bPrLw3WCdFJ
GlD67E2frVpwP2hw8gh9+9vus0A878D5SgqGlB6TySpFlDnDkVvGnscOJkrGtpSuUXqJx49oVWWb
7V8OB7eyiQ984XpMTYEiwEB8L3X1nvvdiFQUteuDUCan1bVnd6HOd9gUrjVgBS0wKH+sSdhZ0xkc
/PzMhp6PlWIxEXNYbuVNiLAhAp9YvDYH8qeZi3nWv+RleS9bUtS2GSNVC1CZdoFfZo0p0wa9r1xi
4kU57D7aNwQdAAAo98s20UUaR99ee9Nq3Z+5yUVn76TR3vqkc0EYE+qMZXPkKvqTqm06GOv86wXX
JmeymXzesUchE9YXSjeZZkMsr+DqWBCBNC13VqRyhxzxbLCveA/WfYsBtHb/ceGqEXkuJ/kfcy/E
bpTLweSCe2S91B2NIQMf9TGBkKLybNRy/kHUMyvuKz9ki332tT5C30/eT8EsAYNUci5tJ1AwWwuG
s8u25yXF2oinayNdOe6RepEBAU7QYqlCzsiKpjVvct/NRB6jZ7937ek/OyZrBly6U2pP0Nt6X0ms
J9+DcqBXijxi5ToCSDp0RfV+hQ5Z0CmnohC+2r8ffCx7qHSSXsOQWq0giQ1tPCH8oiKV6YlXPhtI
lnjaA5tsn8ZNr3Y9x09aXd0G5ClC4HtwgREvvczBWE3VH+lw0jn7S45EhutjOC5iSu/szd6/N7C1
IFUBcMj8CnyuIwgeY58mOHcKu49ly5A10wkg2vfefh5IYLuy+WUxPp/40z8vKnGwgqlKhTX1SN1A
sEaWC0FKv6x4Ak70ysL48AF5azhL5qZdWlRlcOYCyDjB/g/a1UXIZfbp2BsKyslQ20fuPltgsPLU
4RhjKScfOQ7nxmnrMK0SBMVqfohSTl3O7dv/oqh9yJUunhIBLKu1J0AXxbiMd54+Tx+030bJuH/O
DqEHsYYPlQv4KkfN2nAPjEV8qJcm6P4FaYVfixW77K9cgE3AWXjXQ0mc3DGTBQ50YRKNU8yGdtWY
0SqUZt5rBIs+0sRfu3TZe6y1WjSIpg79L3YA43YA3MlxUD6Un82cCbO7x41t4VMRHAJylLfUETLF
X3VrpIyC22IVSzzdIp/0endhJ4VcAZnpYnht7xLQOXqLueBFoFm8cUh9j3cik58J1CE9osOMwnJR
WKUXUw9E/nq5ZmgeW9fIS997y+XLqVMbJ7m5yeRh+cPyf+RwQyerX4e2qAlIVvJW8Z1BjCiLQ7fx
sQdNcnFgRLyd/z+FrJF+VIWbmKwTH6Yuz+8dyxnXF0xQJDkQw1shXbfMz9lFIlxdKzta0Msy8vQR
MpAr3wWJfyoXXg4Gah4geoxhhWiKsYDuWfgy+cC6jG0HfDgBoW0rAVNIX0hVsQrhs0pP6THP+Z6F
jQUv0OqFSzlU+FMCGZ5svmSc47HXg9xxbPjlGgTp7jw6PalQSqy5v+x1CutndFRKlAdsiHFrdziW
Mr9Wz77FKIumwKdD2bFBIcSmYQWaPcbFhoj9UyO/tc70JmG5K7qaR4PpeKu5KJ+VtRxey13r9OPt
7ghHxOSM9TUiPSFtEAmsRweaWIxHDC0EwzRWcWLZv9XfKFzLjYhAmwC59vZHMigbe/jXQ7EdYinD
G1WVvw89haUE2YQhhpPcM01K8iGczfeVr7TtVDjGm7YKe74FCGXgmUDBdoY4x0t7+vO0lnXOfGg/
WR0pSN/AcBErVbKZHU+un+9XC9fTXX+UFYWtRSmNUzkYszBwUP9cF1+cjDPpjFTlsYjtxIubvsgh
D54B4BWlCBpXpkamORNS4u+AOOqYf+mLIsHb55jmqUSK8FBT+zTIGD7k99swj+D2YTg4K01yZCyO
4FSLgF6JjZkrInkgqqqCg1+mPA5CAmmF4wwQWby6ayjNA5ToCyexOa72Xw/7U4V3nF7tr2bU/jlC
bNMAUOVNzRi6Q4CoMCztcCXnBzoF2apQOuS60WvqoemneCgbWqial3DOW8Lgtez+tMBlzlLgJOse
Ae4K8rdCx8iYyP1A2bdUGfi+IRjrQe+Rr1pJ3W0yoexOdlZbePLs5YFiMsOiIcACS+UxyRGQUVwJ
f+NZ8f2vJ9e3++PQMvL/Mc3Bq/DU9yRxCe7eqpN2jvXnP3kKoCMVd7KENyrc2j033/DJzohKJXUE
vM472lWeg8irG/u/XmccWQlpM2vNQdAnzPNbZ8d+3YCveavV62rmPt0dynRGEIOe8e6zn3qVWFVs
638CUs3ZPIASD9mEV3VKFdssB2D9qdXHDrRdm9qjGqx0hFB/9a6gfocR7YIZAXhiJtT1RCKLP7EV
RvFA4vssER5pOXRCfPmU/o1QFfTeBRaTl2evxNaa6qU4/PNVDvIX179V7eTfgKgwUdhGcceFktHQ
Ii1E3Il8+BSEe5nHOA8vkkp0xC2QRzTQl61mCBb1+HHnvx+QjXF5UmWcmUz0nj6NVpY9BdIArggB
ot9DupB/5GpSrrxeRVVw0AALbY0ZM30z6BLZwPsVRzAYuzUTOBX5NA3UBhTc3ZcAkREvz/5RvN6B
YEJmWVk43bfEg5GM9rDhVqYICfudxvEn286KFyJxmqQ7jxXe0UqJbos4lMZzecfHxQAmHtMwybi3
JeIyXQip6BSf6mYKLpwWSEVoHeTf7jn5Sm4n+o5dMJIY2U0uERY/F7HZ181R1CeTlFfpISSashqp
JoXo8d3oJ8rTyBXH3DD2AFmpAGYbqwNHUBIZYIwQ4/0PIfpJNtSzKpQW7YhL/PlIHtxyxCOA/0q0
KduLCpZnO0scjFEcRFatWQi21yMlgmMVPb5yoLClPBlEIsNxSsoyE6ma/7x34fbApbo1zaIQjwXX
7/+nsn5+eiiWn8Yf09q9VH2V3JyAgqbdU0Hqbk3YCoC/3XBhSYjeQkrz7gWMnLqWLkFYNbuRbNFJ
57v98ZnY+gmlF8k7LCTN9wNAugkyU80wOkIoUEWUFQbDdMk3uI0PDIM+Ih3jvzhy3imWx4eqmCne
+5A2UzrVUOODBhem8hE5qOgK7kXAsuYxtyRbXyywK2LXmyLenzDeY/BJzrx+q4FDe3ExI5Xq4en2
lWfLvA1txw9lqcw8QQ36l5AAQ+EhNgmUhYGfkfi2zmEeTmJof4CFt9B2XxWbTfT3xM7gAhjy5wMC
wyGsrVK8tcvwV6EzA4fHMX+J5z0fRHG9bXG7ha4QA9nD+Bh3dobIXNaJ0ZYHCDCR7WBQsHZZHDvU
4bKmn05WtCu29WMWASaZppvyvjzaqG/oR7T6K5vIGes78vHyUohTfdjvnxjLtg5pSZSMCuBKceHm
TTOJV3VKqUOQHrFD9PH8xbbDPFa+HntctTFbtRiofEnIfQdFqf9gBpn9/Cx8ORBTEeotB/+deuWE
RL8XNqRfSkGQ0DRiBtnPLdts/MVe8w5asie1ZrUOps+4wD1lkgu/pU+AyP7AMIoWAy/zXrD6LBYp
GejfzX8YAZNaczgZWfSXsLrPJzGWNEmxRUv/E+tFmizyAcdkk2oIbsd6j+HySfrMRQ8HTtNz/vZm
jLWmQQnaXGzo6nm3ns17QiTGmCmUw/V8BJ7Jv2a07q+4WmhdszMdjmuDAFWkTq/ln56v4qA5IPWC
9dkyvU2pB7cSKAZmfNe47aXA3gLlYt++wqYkCW0TTeGwv/xp0RfDpX6rvEIQ0kzk6Wbq6ogApE/q
tkRuWgF9ibBXsFcTtPE1b86IVDG5C1rEDxsvY/X3Mm1XhKTgtWcF1gubKfIUuzuUUKn30kn6zkZy
iKymij2wvzWSRJPuv30ANmLcmxMJ8HbYKxu/SYwop340KLWpVACe3etpHVCS3ETYYNOtvYaDdpP8
RBHEiIzjTBdanUeJB+pAizjJ8zocgNhlIegXP/4r/kkx04S1tLVHhW7iOET5OjSbag9eaf1fnn51
gB+zF1XGmk0WPG8xPwgQbMeiFsv5PhpDGiNtL0z5WpT5ZMxPuToOnYPUVd7Cg+7UIYNK3frCUxez
hLelV9uw52j54GtIAlr4UZvZXOuA2Om8tINstwTYnxIjQHZLl7F6rVfuuv2p1K6RaVcoJlrx8dpT
uYW3rzGLSwE0SVV0pKAtQ/tTQj4ZHjKlPwpEEqrquIVsU3XX5dOCX5lD1TRxWLd2VBsxhhdFSdEP
ztbqhbnw7xDCCZtI2xs9UScEmDjPqAfaLdmnn874s7Q/JZnis0ROWhATmRwqqBkM5Em+ABYibtq/
AxXFHrhfBVFl/m7d2wFCVVB25DmHQUU+1yiLuIkhWHS3hq3cfs3sdwUgEH983clxwumwhkBivGLz
ijuG3/ufbE70xqmvPAvDXML/Of5J3k2wJ22Fxt/KYKn+pKfzhHCas6tBX7fD5CjX5LIotPM9Ec5A
8md1Y62i9Vvv2V/0TeRKP1V/w4cBWb4TBEyBiOpGMmuFY+oW0TPkUJI08YBhEvOerHgvrhtAY8Ka
jQrEQGo8XGMEi66wUvnnJJUZ4JA0cy6+WjlqB4LLFdNNNGjBXGkl7ofCdQB7DAIEogxpkRhbfoE2
Dcd8nwrICCYVl6nQR+Yz3X2YePd1pTaNnGwoVzgAOBnGtZWZSz/aZstQJQrLyuucSmAoqV0LqjG4
Z2CznRQN0BjwhfxOTALkDG/u5vFm7NFv9+UJV9FORRdSbMrRRLLsxL8hkbZ0EM9Kh0pUXjmqE/fa
cEewWS84bJX7CJfQW17fSvguhFAwhI6zsmisP9VX+ta06Hi9lNMT83q750n0kdzwflDtc6EugEqG
3ZMaqXZRb9h2Iu0kfj47N1+KFp+XRrb64oVmYF2se74bmz8AhGoq+JdmUqBrqq8s8xfjW0jzJ98O
UUyYvBokbgysaNsQKk//vYKZTgV6eoa9zVZBQ4MPAddF54yQel/dj9MWL68zsjBEXFfuhJPY4EWA
pArOuI3FVIKDgow7MYAtyEDIwTrxwitbAdTdcJw9thHAek4PKloef+zFDWWIEdsZNxbWxO/zw7zj
mWt9JVNvC1nHnAOSto2zGZUo3nbgRMcniNV7LQoudRcI7f6/QeETdvfp9YFIk7SGF1hwrceFZLpf
I0y/uDXi9bdNiphLo83Rt44fsfZXGM07pkqYmQGMUqYp1WX7TJ20Ash/LLWJSpFAq/3HfkAG/6i9
Yic1BRIytxP0+703mTQbpWMUY9xd6hbrXl7bmO6pVdatrOj4BquJL2zt4BxPNWwJkAKQhmX68yq7
zFMMvAA9BN5kGV8ks8bjMD5aXYwHr1g4TJYuy9iEK6yMmA19gM63qNZicismyE9y2wQR+AFVHGCF
iCGFXwHYinuUc0jjBgTP3DJSzNUrx0Cpd/9R0zhfNAZxV0+Wo7N81IDvNgZI7fUUISZjM5UE7F3h
1f0Zz/1mhomB9zYbhqpQ8pSSY16SQbbJYBFwep0c7FaF5uljSFlbYZ0/WmHntlt4SOlVFAJ9OzYo
63EY6naHdZNwH1FlmZisDc5UPJUOELv+iZXJE9vzs9I6ihN20l4UNM+bfbN0i9aupc2Sj3NEPvIN
lhZIE8VVpazMwHxCiy/Be2B3DPiSP2mZ82cmrFRt9Y9HyPxBjFw5wtFnlGZQil6ZBvLkVpR03cgi
fjsA+syP2dLijhg7mXr/Sd2PE+kuI9xbodrUX1gQeSKazh2dB3r+2LBoEYBhpQPSSgLHvvK8Bmow
k4jaTGPJ6m9WsNjC1MKye74+b39jHXJmbLvm1gwmglWyjriVS7hgBh1xAxNVwkxEwcIhpG3QN2CI
o6n+qMj5wZE0nDwcYVoI3POFm6wJOxMjY12J17rxdIuhdvOAHLgpfW+f/o2dClugKg0yA3jtECNh
WWK5buULXNs8+LlkYaQALh4aG1JkkACQPb1ZrztBzXuh6akjS1oNXanGOm+Z6lYI8w6Lq5VbDU2X
Bp/jrE6bqgPQmgdsvd0Kru+kNP00FdvvSmX+ZArYs9giB7EULj8zKw/9Z5Pu75unBTmmESTZlk5i
ZtV/Sif67/0qjQHc/D1QuJjj1fbawOFzmDGewjrsMsGxRQm6wclJ83PoLNKE5uoRgL5Qlch/42zv
dciBZwGxdb3SIUqjCeJEyJ20qpjj+HjDfuzs034XEEyrFNYb4FCjEzjlK4VmJz4uVncoZ/IAIDh+
VJ8XjP4oSzgm1mu4H4Jku0Eq6gV8TXRO0pg0jXw5Vh4sbT3GI5z/YYKX26ElyMcKQkrNHsqV4mEi
ygae8s7km+gKPKsNfc1RnqI+CnVzuz56dGgwwnRvvwIwtHt2i/BtCXYFVx7bWsCEP1+/RuszSAzw
tHv0XDMTar81sZDb3We8JIKa04i6t0oppVN6bNFIeNtECFrskTf/U7nJ2+WT8BNyu2OmF6lrP/Ax
JRkRtNWNhMmxJHzlWdlUJoyjTguRU/NBBJMO4gfOZnA1pjU/WQPGG3vXYrC7gr+wuKyrNI0LTnrN
FGHvp5GKuMn/oLtNxytaQJN4TvqMyeOh9JSyObBhsbxl1H4oScIMfB0zmM3HFSAntro+OfhpOJL2
TsIICQl9RN36JJqtOVUsvOBjt5I9JBhnjgAR8W76kzuzHCIwv/e/z+ZX23DyA6J8bOoHbYdX1qnp
uC3dSa/6nM4acxSB/Kz/OpZRewhxVwghEC0/wWvZcrPS/b0vehB4wGRlCgzegqmmFZ79jwj7xijk
RPaC7A0uoeTsopBBRyP9ssN3NIFPTxsllrfPwSXj9BxLZUb+rtSB40swDM41jxMtuQU85Sh+U7KS
HnM4+5Qq4JZO1YjnaFYS/Xm5sGDibguxtXPR7hndD7oWgGR5yOgx1LyemYm9DSrNC3r00PMVwhrU
M990/okMb3+fHHxdQfwXB8DiygpWJkcebVRhbSC4vFKblxMxah0F62f4DOC3Rp0n8P4W9LXtdhl5
1ANHFyvybLjvrzxSfCLe/490JkXN7TQkNSrdagJ4f3IdPdOibIGXlhdpGi8biDG3g0BQIPusZl6r
XNZlHUqD2wmZwgjsqh5W+ml5oRfVHhELj90hdC3Q/GEXCay+vVVcbHwJXNwb+rMe7R/CxcuXVIZB
tRm49+A8TCB6RejzvFJVdmqZB85dQapQxUGVGGjx3+X8WNUnyeAII1S1zwZOueTtRKRm4YG7XZ1I
RH3XCQIUo5CSrkXC58LCmsm8DfFAQpuZ/IxAsWl5+zGn0HHg/1mX09vqUbAvpmtOYMnWcFFFuIuh
8mZMHo1/yn1IXknqOYqmowiFbjLKPsANMLkkGQjGQ9FBz/5VKc4AFWUXSsFw6FTHzfJT9BQIEUd9
3DCFPDOWchUB2+sVPo981e21O6LC7lHc6qw9uZXruCgBLL+5FaiO2owZtDQ5um+t6ySlK74cCRaj
+d3aMa5W1MvE4PsIqAszFBiwK2Xnrhr3fRryVzT2sJs5QN3Eu6YL+f4cjn+cPwIMF7+t5LX2T8X4
kUbZxzT7kElYtCi8uMPMfUuZatVqRwVbWuDHjLZAAF9fD83IR4rYQXgq/zc3Xar7wEmUXxB4EMUI
cpYh2UPRCXG1akPbYH3WmA13mx+whJYFFf4I/fazXdhDHll6qLoqqX+0J1qDWg9GW21lpZTWNRAZ
EwXAdU2PexYqSrXt26SyN5w3g4ZNh8iakWE3TfUYDR0lyIMAdWj4otZECFE4Szn7xGafhiJgQbeL
vL4Brj2eEdrtSNiesCFANYhRYP8Z8/QQydnDLJh3ohqzYH3oUZEcg8UDft3vCNXwlcLRwduFHBW9
7GDEnYt/1tta1vCoXlpjNtzJtjD2VsRjne1L5bh4GbJ3JOqaGdF4wpW/fNnHn/4b6NvWuM6DAKqy
UzqLxEWiWxcMX+K7sbdtUPThcmvKnqfduZJzkiozI5Lpx3+JfZt7mCe0hYOuST7Xjo3e3dIG/Vgj
V09d9cz5i8B01JKN1NgAEgPke03NvsNbgDzxB+f9ZKKpaBIQ4sYsE/NMopYqH42bpNwVv4lnx8/d
/H3pxqcFBg01+R7HdUGtc/7mVyqvV3pyJseMvcDaL7UJp/9RokHm3Bmi+sDr+28rQkEZTpTZQpgn
ee8Ug0VmdK3d1CCsKNKf0ozmYdKdKfP/5sSaNl/QOE8ifY0rxcvlCj7hWmYGBtVXuXvooK/byIlq
E7iFIUTL4Be8skHVaJghxMDInlJxFPFLlp25DO9uEyXRS4BAOEMDWG+icThLflRob+po0qDHwBay
Vhjm2O6Ef00h7mNYpJt5uNqhmeCicbau6GWxnkE0LGi79GsP0L4HJY1YC+hsFRqvO8Cda5L+JOb2
9ZOSLS+V8wR3iHcGMbW/oXE4NGBHeJ0z11qL+kGfgYCykO/U8nckO6NChTsRs0/qYgtAtnPXaLvf
C6CgqLgLKgxsQMCc/LzJur8KLGP7pMCADAYJkwx2XtV3M5DVUIZqdDBmPIu+jGmSwySZ774+RJFH
F+DEIzcVWgL2D9a2YGwcoZOvUDzySyikbTXkZrk8EGLNA49HM0JkdRCTMPKZGlXHXc0rJtarNK7p
2WMIbiE1Fvq6hPhBN3HYzpDgcKB/Ur60t7hTFOf70WbZiaExQaTHpb9hPGNdJG7vUGFgL5UleWV6
DDPIyCgsolvk6TA7k4QRzUxQ7i1UUiw+Yag44QfbNwR2GZsCeg8p+EZEIXcAktdiowGG8lvJaEGG
Uiy+fL/PujdZRCvVxS/JNUjylLKxv/LpVd/XDCcaSbiOmoS43w1IYgQM4yRP0zU5v5THN2/u8D41
3N+sQoH3r8VoT1QXYNdQs/UhzIX9O1BHXsLVE8y1mSXYX5mw+LwY6zIxtpOGpFZTXiTkEpgIfl++
dI4T/Ke6u5Quk46YMArYzL7qLdefi75MpSZc756hmLle2JoPUhJNAtQTp0fsJt4JHBSIrSd48e+G
V6IiDX67F+cSgfFTLbk/xbtjc678fMEXOiUtXrnJ7k4Lkkah2/HLfJMb4ZKXBzh7ExikQd/fCShZ
RwE8dMBqgNlItbKAQorTupaFLkli7IvJmk1QZ+YiCmdtpI+eYlaTnqKKz5M2OuOimcG8lZXjgPt2
T6Icvd1jJQS4n/iyfa0/BzlWEe+ACOi300GdTFsFD2LMBTvpuRNbicK202uaf4fzQIsQxL7rU954
4Afsh36hnipcGERxYnKdXD46DK7lboydNX39ucFbakteJ0ZhUvR12fOpFjYsInOk0J19RsijRAKt
CZtJeCmcoHHT+0Sj0m9ccPE+MP7a7oPZia6SXbBxmM5F4PkwH4EDj/9iLfGA+oSBXe8ntgzNiDui
wO158rDJ2neavV5UjKoUa7uRp3NqRznpKRIHtlEu5bkYq/i5mnmjAFTShRpI58gDZ2ETGAEIYxkD
pVyFNu2VMe5d1U3IdsgLqQn37C/ep73EpETi5BLfcMpoHSCUZW3wjMTMtkNIwT5/VhMW66UaonTJ
JGXSYrDHFJlO2fDL3JmeSqzykjgXtL7e47NCH0gyro9RWrU/+kZmrH2xfVqBrNVCcmAOyiyj8bG/
fGYICnh5EaQgTSNlSUL4b9aVywdf+4A6e637IeeJ5TUxacPdV9BwbCffQf+LVyO/mk3cc90u4LUc
wMbkIQLIzettZvuJ4h7LNMNjaOwP/zfqd7PgQ8FTLqRkJrBAI/cGtP91BMZGKIKYxFr3ylxqAsvY
PRE/VD9KUs0H/ycOTe9NpSbTneA8lB84/LTgnMPUmpVW2WTQGEykY+4HA5VFpMvh6rdegQ7WCf6W
jrHqJezPPwqsnp8rEl4h1aSJOcEWrN62ZJJx1eW+JkvqiNdQS5vkV5pInbLo1RHnzJGZ8nkP2VsV
2MjXgVsbX3rc37MoJw6R5Ac1JtwvEo0aRI3dgD8/PDwezLvkpDPhs3ysuNrSekrGXROa9cCADipt
uSlLyVRDecFpmfk37z19ukZif/Hb8xeaTZ5rhKKON4O6i/zQ/mTP1SDRjO82n7yHn/0+fqVLlC6q
rBBu37gt2oPeNibPAOYJgmrU/Hc1kvMWIZjMvKkZtGvgFktokKD9C2FCTlAQuFicpJQKPs5EI795
BrYCVi2fGHTHM5+VbXDEW7W7yoMa8j7x/xmmg5niStS3sHbCn8pf9KxiapoQdm2LDC5LYZm3j9Fz
lZ93XQ+OT0ZG8rTX2f3GCSkhfVlH5j74nVo3vkVjZRHtJTcWjHAq7nPSmaWIO7X1BiEq7u0S7La4
t/AVSmBZHXEjx5fTdV8AT0wOfQOBPOXGS0S3mB/hajmpQtALjF1KFI9eX4oUsaznNlBjyIjykoSd
WcAglP96HuBS5ZlWuVV4t2j5UtJgESPG4aL1wmqKuKfAtedJ+6r4o2HT/TJx8RXV9eMrjVAoGCaE
l7jyTpoKL+gXKumGNIXTI9ds+/50V1dwg0JkEWgaWJbr1bUlkOFK6SsRhU1cXLKhwyBjBw0QBlF0
6kcsWDLC19TIbysPAAYmaA8zqGHZnvOH/0pQQsRPcq4pIjekomYCCdP9yM7bqZglQ/IhRCapuJFG
wcVGbC35DFW5BxOGzFTbAA3gg2es7G+BapOpZcZhpGZEnDH6RfrtN1N8VUWw8kHbu/u6/igmAXcG
EEmZBroydz00kYo5WENimgOQeP7YTwAgIxdiMNJLvI0Ney+AjnOlcZJzLkcn6dAjzCRub8ro+0nb
4XElCOM3sCeX5DA9jvGzqNHE9OlSnTZ7g6Jz8P4k12u59oG+tBdy6ZxElrNkv9mC4QlyJC0N/pBE
EDJhw84VlamFX4UdBH3OpequDLOmKDgHgmCQSkeQI7repO8jWhkyKhmDiLZyafa7d9EY4JhziDi/
VJva48X2T8abiqC0MsQvZWqeAYfRUUg9qdIz5IEzRF93ehyXjED6+C8O1tCJvPH7ml6NTvZh33yK
b6UTh5eDXbD0Nrb/IjfPsVYsFvneaVQ+ImQes3hzrG9ZlNZXOyh/ZTYPTwecjJC0OurCkqnUdboW
KrXSIRRZO1/0b5VvHpDkxVFOcENBTgGe7uuRICwHzBVZRgPCqYVgiWRbPti/0NfEIadmq5k/tOt+
lpqHJTHnkUzlwjy3zRQ3H5M1KBXot2Yenn/ok5M4WNlI/Dha0ioZoIWkFz913u/90OO2QkraSXAg
uXzEmF7dnhUxl80G8pOFpDdDTMYUvU9KUP4414MXQhIrlKS5K4IBghLbfekZgk0hAUa/hZV0YhUV
gO6tfQoiT2V6JfuXwJHWR/hF08TMV89DvpMgyQfVfryUO9AOR8CX/jjvp3MI0pGVb4KsH2YpDxYp
+TkC5er04RsOnDUuQxOXSsrpYY2H6qMdAZFGLdQIOJAJw7JJLiujIhpXbUua2nh5kyhWj6itJNSH
fJOna1ZGCgoPtIlxhqPI2qHoiiTPfxAzadLnk8am8h73W8Jh0JtPQE1BxVM/DZGiRIs/qjseziwH
qnv+Q7xkgeW7xISd0SCzSd/7CxGYOYMJ4cwiPupvXgT6p8fdV4O8ZCAPCrVeEq1YJkF0FmVbO0Kf
0XA+3QSQ4+otEE3dUUe7UETDLX4+FjAZjNoYUlQANOCqFqAhGAcANOtzBMcNZg9sbWTvWgdy/Xnf
ukNreXDLtn6AJpYq08WKYCRv4n5on+WhSv+X/BZ6AUhP/5eoCjLHqo8EhCCW99xgycXW1Fo2/Uje
ZwqunLWXCNbz+Iea9IemLfCerqFO0h981vkuHT7wRUdJ+FKFDoNonNvTeF3GmoFPvwbCvnTdQMeS
VYLMqDu1F0lCiPMbYNB9Ktf9VDCoALaTvyHLB4gwvU6oWuZ/RUN2Oln42VVClKshopfOU37Z24+q
ika5Jgkvdf1MbN9waifZHNTcOZfDaO5NNPFGcvMo0G0X2qwm1/sK6A6BtudbsUkprzP2dhVq5OP8
SUekrr0HBxtqZEhrOC1o7TD/vUBpXGPA/61BJ1MdCNnGiiaAxOYdSIQJyLoaQFf27S7rVgFzRUWi
isDioJob68mYyOD5Ehog46iGFKxa4TpvmcDTFYB3O59gHxB1BRC89GHbmVqDtX+pzjsFzkXTgzti
DVjHXakoI1D/DbZwP261ViNNPuv1h0q9Y6OCXm8PmbMKKfoz0cACXyTm9ADBpS+vETNnFIm0Wll8
5+8cN05FDUFK2PDR/+l3gvjx18WALcGCXjCxVGxRaNiLP0hqBg68McpM093A9yqwKSsI+bTYPCdb
gJ5i+8DjR6l05qagE8nypS7ihNAyFNAQR/4xpEw9YYgRN8k83mOUP/MyP04bp/bHpsLV3VlV1WyM
FrHbqkSLg4Wv8zczihv9UJSDDF1XbI8c+teVQ9T0nk+cB20XAtJpEDKKw9iU5u+AS4WtDoas+Ge4
PKOp9OCyvOz3ODWU0zs30lFcs/p11kRhBTV3nBJBTSbMpI9L/HWfHYEaxMcm5AZjDpzg8iBfFhZN
v+ZvQTwlPASx+EL75eZv/DHCypZxonujUNtc8lJYZHZtiFPfbUSKWOaFoG7DLKy2MVNGrTH4ZvNk
zhPnZOTinvGfNVL0e7ME/1DSxiwGt8NlzswYQ5t5cbkAqH3VxsxAyQi3/gxZLAJ9MLHLCxIEOmnp
dqu0Ff271sWWWeqP8+HKHdhEKwN/rIxQhrZ0/lEfLyJDxDcV/3iPd3R5SQpscbxgyG5bQ47D4aGV
/S3aDyf16bR2X+KPbls7CKYou2KMTh5z+3HqUwoqLQ5tk8r46eN5H6VZlDSfyJFrNltzTtBe0lMZ
EKT94t3BZGtHpsZfaYoKXuKNvLiOywYK6kd0hfB4wD/lqkdRBcQJ4MMP82BfMXu5Xii0dn55IKtT
k0//TTQ2pXlmXD5X3m7EgOLH7dHcAV/p9aMlvWvfHLVprhAvXuF4ll64Qoqv1ezo9/Bf0LGaFBh3
MS83X+UK1lZF1XKhb6YqFCScgFn/53KqE3VnmT7T/ihyQQdMeZZJrZg0jkhieGderr15Zo25C18E
4v6RGGvvUno8cYI5SqNF69iTiCYuqQHTfYmGcYLVancCno3V2bXvs3Px2JpahNJ6iuzS7qqc3d9s
dvKgD8CGZ+j0mi4Y05/lPDgPb3hSlqlOPfOXq0d/x2qEC0l1dEQ/YnUUwqEoe9el4nmqybHUfhsI
z1rENo7uppgWCty+cAgPDiKUTRvyvKSTxFeJ3yhY0BJ+YJGIfclTQtTlzKetb1fDCpEYdjUycKn2
nqob5PoYOsHmcOnH03+/xFyg3JLM83NHomwKz7abzmbhJN6rnqna4SQgRuuRLD9a0rszrprRzVos
1fqSKfpAnYQUx0P9M7FkZ2GZn+hv5ZgFsOrAedbyUCNCa8paEt5GiYykS1yD2GN+AkLnNqZhhLml
AeXpjZ16N4QzGYSusL6yRLRN5LbpRH6YW1iblcpQMPOCBUZTXXIT9vArxKyvufNnruoU/f0wJept
NRh3uRQYaFzmSxb3GhKdFoPxqwwV7+XmDuQ3tZ217XZ1EwlFqRqJtrvAa4XHPBpaxIEfnDixeQXA
dlOIOAcye1tvuhqUnzeoRFjb+OX0tAmQpHMtLTynb0TuWQc0Vo78+SkwqU4zAPL6bK3F2gyynrkS
oLWmF6twNVH20n5h1IlTYgMFY3BXdxrMa9/ihJnwCgWj0xwK9o5AlnM/mmq0djG/kiM2sFNy0iwa
alwXKtVOXND5MiB/NuASMtRfCMaoLhYSAoFcz509b1sZk8KQuZ7Yv96Uyb2+a+3jGliG9LxAzv8L
e5cX7RHBqbYJ0GGqB+Xd6db3Dl47rJcrpYsPGbGxd4jPhSkTqo2GTzBn/MB+FPf4hcbr+hlxAy81
Pi40doVxI/sm7MKBkJvYtfc+h/6DzW5fYfmrz8ODGl9HWZwMqxs2SDX64G2CZFtzJIfQWigJLRMH
W2usSjqPKKzv5quZpDo5Fk4o0e1+cvkuN5KO1UZOrKJJcS8xwlvITHEalUuoYne4+6LxJkkfGbdS
yF982foClxNpSNQtG9Bgg8SIJmN9jfihp4O43QIoREE13tLspJU52vKEGqvWYyiPwwvAek0e6/mZ
o1qWZZCpPEUNWIxLoAfFmui/MzboaK6UtSV2Nb+1yo1TjbBjB/cwCghWRUZOi8lEerAWoir3EJNk
OI9Rv2j7FU0GVEKl79QURYc6HcxuIZ/6b5fK0s3AqXqS5TtkOHWJppW8GsLZZH/YBzeJ0uue6I5h
I6b47SSOBTAapWzrJJ+2DjcH8AAIL86lta6bV1FVlb/MjqszS6O2fOHCfA8lg4yoYK+rVKazebcu
jTQI8dzcWnqibD38j/2J6xq2MjajUUjWtxtNf/nqokStXRGs2WRgZPm++HWpUJlydvCSYlMDw8FB
4oufRUZBQiafhOxG//mk8dICCgWZB8kpIlXty63ve5EVOY9Q/3XdD+Zg6wwRW7qggGBGQBnq8URw
EoYpxav+0QU9Et/5wTeuIdrbRf4b1PjsT0xDFEeRUUgQgDmtoSm7GhIjd0dBp88sfPqU2YpPkXx0
4thuBEtGy9LLLznNdyvXwPpzhxDJOH+qcZCr9+hpc6p2RM0bJJ1o8Kjoa/YZEvokPF+t6cal9VDX
9YdEXTf8SaM/jW1SsGFFX6S/eTmrxw04OB1twza17EPG6OBoVAjxa9c5gtVrUJyIDC7MAbm8CPAc
4a2rwlGZJ3Pxnb3idkt3pEGWV7n3L/QlQGRE6SrQ6x9CtuyIHJuwzKqGI4lvb7JioUKDMfGoJCYZ
Vp1ubn0+OG8IfWEIur23jrNIo5k1kHTfHJ5QVxdiZdXzUHOogXZl/7ui30h22FyVdCiVECqwf7vP
fc5pIiqZ8dNgWyljVYdvFWC66x+fFmYR2NdxxFMRlTz1AujmW+zvRwiYmxTjwLIIl6yglOQaF9oF
hGng1kdzvSFmb12FO4yfc6c/Y0Oj0SzV6m9z4UvYlmQNDTuV8HT71SkzWT3Dfy0dI8G1WHZeqXm1
cXmG+iEtbugQZfm7nZ6BVvJoHaS59h2D0AWgYLuCKBfdkCdSMFSH0vv3GtoR9psto5l7OhQIo/E3
I8aNrliIkYMaVwaaL5ykrj+26ik9T6xv8VoTBA0VmovO4PuHRoJsL380dDWGbDs9NBP9CAltsRWJ
LIPn7bc6Q/SDUzI8NFOZU8Cbt8xusCzsSEF4GvtXSPKuzYM5QAnHh00aiNO+MeP4xnojNDBg3t3O
BNBUVWQlf+jqyA26vZOrgvt/Q65xzEM+o6dobPL+awGGwHWP8fUZb0dutkoxLyckLYcsGmJITDH8
su4jplrSafLNlyU0S825XmfC2XcYzDcDB6uoRBsb/AHO/hXMNt77+YRI5tT/Qyzci/dxUQGL6Ji8
XgKyRPo8EdAvFsVH92YqS5xIcPmo6mUElOh+/hDzK8QjeU3Q5+wyzBtVHLL6J3Cr1Z4mAxSUyRNX
kodWm1IvJsEispuerRVHN+hI7WZ1yvZjlfU8R+/SbW+xIssWWHkub7E5sWS5Zzq3AyXH3LPFDbbQ
5onVb/K3DN16bOb0H6wm0e43teDOUAWPiYVEWSqzBpglwV4xjwiWixHmuBPtQn8OJWsueNKgNi5x
WfbLmZfscpE87yajaODJbv300H4SLFSYC9H9xfTf1+Emlol9izEJA8YIYD46K8EGL4JVrCoiGMZa
F5vqIgGKcOOgS/jeh9SPNnxQSsbpMGly4eI7MvZMfPw8de2pqH34hDR7TD30oo9Dv11u5Lo8zTQk
svhNTBJa2Goe9MBdsbS4aTvN6RjxZkwRf8u9LY58efpnzcKkMaog+5FpwcKYNpJpnlclkpRrQ1wM
j4w9dNcETUm8GMvy9h9s2/oo94XhZQboWDq557my6+cQqjxyVzpZjxUi4iXtrw8GBn7MG+BObj/Q
UBMSE18cH39gp9/zilWXVtEYQw7x+Fbm3iXLkGaIdt3fQ0ft9o2aFEL24yT2/dv0ZEUvEoJeDytl
gwPxYt8tdzj56ea5A/Snc3nEuNwXorrl45qKmMfVeuUX5ejT2qgwdqsn+IwSOAFlSrYoFqLEbQ2m
Lum9sdZBTLBThb/m9GVbIhfIP85LQoAthMuBupwBesIM55ha1y11ssLixzETbGbgrkG6842+IxU6
Ntx9q67UH4+ZeMcLwjXBmXlBC6z0rSoLjOpzS3yrc8xy5slHerIoyVS3/rWbvcZq/+Eih4pyRoct
aZrsAFBxGDoZEmXmE6FvfSAbp6oPr+5Nczc4aqsUNApYiOFKj6FSlF0B7lUmckkhFpTfe0/9xyfc
vMH7o8+fkNvXaSPcviplxOVzGwpZMLgcfUZsuKyHhCUyGQO4MH/D9CgyVQciSRBNm9MmaMqwn+3f
6mQw945Z3TfTSk9wonE6aTDI2dNSfTEalMvahptI/qmPQhgyeKWfPfrduD9Zaw11Efoo1PbkfTFh
C4vzgU10gQbwdg/nebC2GKxLsxFGIHa3KViANQh2zqxKTdwRlVfMQ2y8q6KwMHxhllczy0Pwm08I
YDFWac8/hk2bv6EOkHfvlZHeyNHKXobRKinsloBbD4Be8kF7MILLqCSWgdAxmhgJPhK97oRYKPLY
UEJJyAVUySNUMENnOAZQRy5tC+CUyiMb4LSnl4/MKucXZbavp2sj6938ghnyhx29Xe8MHFQ12xS3
vAZVA8pmncpao4EBl3Ojsn1dENHAVFvwolVypLdyXUWZqqSNuOYZwjihafM16pXlhs7KaUAv3auM
DhdFlmot895hjwgyoHLCH2X0ueFFu9RF7D0JV9QLHhW0bbU+ooR388sPZCJuuoa7TO6DtOEaeLgR
Gy9UCZ0GB2/HQih30sgfVcghxwJ/J5XMJM32Pa97vE2gflbiQBAY4EVO53Ni9cWHX5c6C+L3m//W
j9nrbq3J28Q45D1z5ENvAyW4d/yCssVJxh0WmaKv9LdiWKrr1n3NkuFovl6S/1fpqnd6icUXZnkO
znBvFUD2Hcfl/6h+PWGKIBQlgWHTdjZp5ZDylnGu+O086z3vpghxIG86SQIfF4dMaPd8mHDkbA7g
1XHdHCz9yLjjBHURPBSpXmaRoa47DAAiU2MR53cRcVa0jA0+pvBkVBnTGBss7+c5WCBD8uIBC/1J
pGvC5Kqm5o+MPJaavXpATrLVgNyoKsUCryNoW3WLB3mQvuB8UtfOMv0vz1mPPMk1Y/uEZ30zDx5T
jXx3y2sbmdqclF/IYd7pdNuFrC6kOH+pXyU1/gs3JB8xHNWco8wdo82xvbxBsUhs767TPkxNdsMh
837+aF6DnYNCidSVxpijJPmC82ToXFe9Ez+ud7Bvli6biQIjxLI1kqPmYUDLibNPEd6TL91QJ8/4
U4xh+JCtC7axunhE/ikYllwkIXg84vfgJcUqTT8crbmhd9NtU/UNMYfYEm+nzrpF9XE4b8/7ntFm
cQf6UunAbxu8IuLKnRflXMlv17iQK0QcjMlvpe+xF/83KSTnO/t6zCSTYtSjI7/1xxisHXc03EE8
0nlGbCg+OwzGyzllOhhPQoN6kY40mxDiqu7Hinvog3Nt9cCrYjTK00LVzJWg0MFLygh2uGcoNm6N
TPLOtQrd6yMgMqK52FKrEqvZiqU9EtNVAbZ5nZxo2SWkqTrC1qHE/m04s1/KGNc86zHhEqXTXEgr
WR9//flvRHMilWUSYF/2s/gJGMqKXFryKINIn9GNm0Scg63vXHirf6iGmeO19ao0VUwsOwsEYPGo
x3stmVidP4tlvZPypVVmKwRa7yaWE7d5xFa3HH0TWvvzjk8YQCPT9VrkObqFUUh1tH9aCWdCSSeT
Lp7Tm7AO7j/0mh7nJ4aGvFJ5lxMHXu3GhlT/rIIphZV9z+oz/6fdwgAssrrKFYVgX+vocKTC6Hrm
Bn8H9mD2LuoSMglhEcgGvE7c508BlpDqpFgSaSu6WM+dpgfNLwVotiHRrEQlMqJzK5Vsbc4voiml
RX5aEPa9JcFc0lQwfQoB6XMM9wvVzr0k/oDEX+ioAwC5My55E+4aw63W2FZPU4EYV8UEiq0ZeWlp
b/yNR9+jt5Y9V0TSi0VeSG7xn2qBVi8BHkNhjpjBGeAbK5Vpes9GB2AyreNsaJQV8nhmRYjpICYE
zYdyDPpPkss1IPvX9uwTBIVIC2AHI6AguNz1xiUUNyM5099i+FIwE0G49Hl1q2BGYpEeSM4PXUep
maIYvHUbgyAsxrSmaJkyk+3O1naCjowK1ZFk2rtkVChuqAgalNevXTqt3oFRq05V3IBFOSl9jPsk
KsX4m7IhEOZgywnOOGIQv/VK8ILL1iO0q1s9EWoRzJ356RU9BThYH+AGCPqJDNkEpsEMkK4Hm51m
nwoN5pX4X+I8cxeJwOnhscWiYqOY5KXVGFA0UlZw+bcmfjXmnYquLt0bimJpv3EWtndELLW9+XBJ
7bJ30aq3WrUkEAxpo0pkaRdmcCQCctqmr8kLsRSxfGbFemwHm8keedysoGttTjsMzFfaEsLWm9Rv
+xUWO+vcC6MZJ5yjc/KFDeYjtua0nqD7Tj5j52q0WH7+Sc3asLhaUzkjw1TzJ9/JnsD/1u3EzaJz
EOh+0tXTuzicw8QESEcd2ZybwAMyFlfH07FVwXcLw6ZhvugJjA3Om6hyEaOAPyzs3kpWjT6kUUac
JwSrjCGgJ8xUic7LpwvQfGigWCDO/oEpLWkIw0DYt/1Lj4D9t2F8KJVNP6bcyTg6cCNRpwhy01nq
02DL2y64ssBaKrM3qC4FseZV2Yr1mPs9IycZgmhIQAEn/I2nVYktH5+/DYqXnjYNFUGi1PIQisOk
de3yOXxqzEVn4pCqpiGSF+ISBTCyE6xdRpM9nQ9ADDjZWq2sj0vrYeX3mmpng0ycQqQVf0L7SW9m
auY3fLxKyUwISDzF5d5wDcKFLrk4VXuWHJi44XgSeLp2A7GOGer8mjDiGBj5F4J+EOgos+54RV+Q
gVsz9ZsZ2pIvkuoiqeiZe+iFpHhoWidzRPxlu8ZU21R9l5aLClWya7fwNzPMisvx78adf2z3xLGC
vUZ1NUVTj8sKRdjd5kzCIXzRKDkFOROkaIZNggyrqPV+36fIz9MpxyJaaiksuvpLGyoufyfW7+Bp
q2yMicuLeBrDIyte0+tiTU/vOeZxIVfAR16k5vW7z8QLB7+sAIaEom1iZVv2UD5SSbsREVmpcSsr
enQ+NCPeDeQJ1jLbmZ1HArG64rqY6jj6AcAGbpUpSvX1ga358FelmV1DpHKS7QMdViAWPIwGoq4T
jPl4PtB7dqeTSwTs2nL+bul5ygP0S4WIGcO2+jOKcBqIhAYc7V1PxgOT3Y28lehXtzlG+l/XxwFi
8Kw8IoeYmk2JaQ7u8w3acgIyIpG49C28usHlOzkuMInExwFtbDahDzVLGCsJldEoz96K91E92pMv
TWNCUT/N7Tb+t5ivI4/CUyhsCjUxgPjPcq/mmBs7N1MlfhmgRye4+Js+IV+I80mb4aXvU5tit+NT
i6QvrJDN2SAsu3ztEE4u/NgXTIVv8AVghhIbdQv6cbPA6WIDij8hkdmxhbVjBkHtCPoVbeJlCPfZ
KEriI/WwbG0HliJcHKJCcxMUp2/kNl1+7BdIb1SA/Qnn75JVxLt69ZrA0Eg2WFRitNKHq7ktzKZC
Ag6CU7w0hyujRhxzwA/ncxJMmwi6uePNlIRoUycVz/PV4hz+ZSp464J8wpbMhfC66ZV/mGm+atW4
AOU+hI9sZVJREOny7C+ROMUcsClWbLTSiDb84ncdrcKUNfo+NPVm4+OoUfjtQ18dbWUijLFAquV/
dg2j0r6CMCs6CxQ0l8Xa7sjolOz1B7Rorr/NYxerdAM0mR4WLleRtk5ghiKNJMaVcJJXzNtUuAhF
9Lp+E0uhpJcwLAFcGOJRB+Ug3dS/uzR3S72YxiVwRenCnHPZNMY3Pqf/m8watDW/CMpbykvZLFdB
O9NzEaZvB62a9q87a7KxRpXlUCOh/fpRUs9o7x+ptxR7gnO9taUdJ4Jn/DBVmERfFmhhytmign+h
v2I4qoWPqe96wq9tbYyF1vNYjhVTRhQZc+NUNYpxVA1ML/JyO3n8iCYs4LaZ/tuNd1CUlQXEgi08
pR7SHWSYVtZ4H4VUAZFneAx5LdMtar2qW7WZqejp59ywkyEH/tOf9qaCs2M72LsIsq7cA+FiFgjh
9F7Rw0lrCzKGbwO4zVrIayVpJdOkBF/I7BKIbJpD1N83v/h9gZPJ1UMBMuOYDdIb4tLk9UG5ZJP8
1GK8W5iQmIeLycYH7VgsycTgMVUseMq0gkLxr+q9+yXuaOG43/cAZag3CMPKfoLv2PzYDM27ti87
ue7fi4GPa72C1CUb/cQyoALC4Rlpe2ngqm/OZ++K2KhKNNFlWl7JJPC/xCK8kQIGZZecaQJN0x5h
jzwOSWXp7Kaxxmab+7soUILETM6YOascfAGGxzjtS7+vHHQebuoOj48cWJ/FlGvRgjjuSfjyjNDF
jm4SSxyBE5uJYB8YalptTFBb8eqwprRjAhFkIJoIYHX+m0GhG2/1wo88cwS6zgRVIVx4RF1xQ055
d5rJXvK+fJZh1V/Z6SbXkVSXj9/SdObpFqa5cQOI/sfJzvs27io7jy8RNBfsGG4pGnKnvxmqY6Af
q52hY75e3dS13vKeSeayWSM9wfx7emcHF7zMf3RfwPMFYAG8ZM8O7+yzinN4fMGo7XxJf3bsD1IV
L/RJiQg9yllnLDwt92xAsBQxeX3EQamuVz+YGoRjxmAcMqkVNL1+CKdaKOOTlTuWXO9cc7ewtfRK
uGFAeP0/BwzObrQK9PE/FY4pmA7qEzWNd3Q++uSPHOgpj+rl0/P5Mumt1afIpCTbZwlO2MohUxHK
K0GsvZbRLGTBo2r0eEwlpP38ckVuBCvpDBL6TDD/D0XtdnV5PsKZq79yegquSjvrABdc2RtydtvV
KVfyopSdBD6cBmSDjbhbEImuCoFTQ4kwt1GEocl1lQ2b7tHQQol6zeL07+sb1L1LD3arnCj1wByh
wMBM7OwZgMeK8BbWBCFhoNJFxQ6ufx13QlFFXvpsg7z5lug+iJJPVg7sbBDC1FMoINahGeJKrCuB
d0kkEZluVVNEprj+kLxles6zKldeg+Xgr1rwZJytMqHGrssPLZ4oCLOF3BfkjpRAH2xuGYvLKKak
JpJm3PTMLSovo5ilK9tdlNCJBb8VlRAZGu3lhkXq2sNPCq9usF6MDKfcAd1C8xkgLUugTYN1bwIE
8ATX79eLe9vCfw+kYa3Te3d4olG0XoSAYFvsecJpH5TyngJlxLXU/jSFNkcSgsWLVJCo4/U+tCeB
h+4ArB3M31GEPfMuc2Cyn/As/ZlWisOqNLwB3sJUvvubfv09fxkKgwfy4oj18YK5EnL5ZzBueA86
K1YtxmywJM95RwVOohufM6t0YqPaaYdU980R9mAorD+/aEoysUPQaiPTj6VYd+e+xI1UvOr3LnFc
Dnh2kCHJzj4uMQhHBunm3ZAITRju5SytohGsyE2ReXQMLTqpoGmo7lfvIfYznSZ/2cdSSVz07b8v
J/672NRASU/Iy8tUhBl7s+rxJ+iTuD5HzC53O+kKwxZ2xjlIJQLaBkWZqmDuK/RS/noKKph4Edkv
0kMMhrPiHIcURq8AZWi3LwQ2CFuP6aGBaknn8qEJMBzfz72u/eIpRSt5JN9qJpp+Nnl1ORByFyAM
H59bPXL9uVSEuW+k0mofBXOGZpuerIqyVoELmSY02UK5qSHStX7tpJ2cBWT+yqr/u6nLp9kGX2rD
ULrZ+2WniEXX5dnDeGvSyBx1MT+jHQyEbAfSJkvWmiKt46Bkk2zTWwu81cHqtnz9rGUeUZXBCOv0
l3ski3Qg5uoaEHYw3QbdV5tZRU9Gw29mOJWEl93IJDcKJev7tr5yJJgl8SGXvpzfSKDQ0eKPFSa0
Fa3HAW7rPwG7yjAUIjOVSNvafbxm7P5eFx45atF9EMLXRENHXoO0lTA+DQiTqN7C5+C6OtgGdbKG
FrG3ewFnfUqX7a3FcpFdpO1QpR+cDUA5EoqV8Nd5rI6wUpwwj2HJfuvC2F/W24x3TTEk9bD3+od+
/3fMkNquAuoV5wWiEIAD3Z6KLoMJOEm40ctljj7aSlTGpgePfwZIu/xDEoXq/8Vma/w7vNC/A5U8
ZfsSvDws7QublbvvQe/8OT6aiTd9f9vfLVYWiz0fHcwAcgsnF6zvVc1xnHx3QUWvXCx7JLdHNxhQ
CUzCyYGWxMOLA9EL2Y3bYHHERVURpxpugijOVebavNz9jjV4c7dT0aKd//MJ28hB9oG/uP/BXdTe
nEie1MS2soTK2cKYIxVI97TwGjyuo1SGlL5nlbWACe2FJaBI8tjGkUsubg1r7dp0R+f1hQK/vVQO
B+SyrznhaoqiC+P8rOB3ZJBvPTeJ2S7cqKc2MH4IvE+NRbgvhTnHUSifWF/ZVS7LRN5t8gVJ+QYz
dqajEB50syXF64+uymdmqGG8NuxcVxltOaqGAiMlRAzKHRmJpWastrUsOt4cRTNpmstzW4XjJn2Z
BfpCrRHH/L/fb7ahDeloITiX9feg9Kg6Ai8CA+7PIoaceWUMjKidTHcHBpkovnpI0R4K1yM+ndef
8/EKI5zBNvYYUp0KvKecDJMRyB9Lv4cvx/mSy2TPRZF5Ah5riMf2DRj+WTWMjdrhsgwLE+HnX06W
UiNiXQkWi3RDB7mtrYWTCq+m1bFTLhYvkrsOndRNwPkhagvioJHjfWJfzykWpbOkGrV07sfJtz6J
//oSGcCRWRT+7WRZ3BhsZQor3UOuFsoa2nKQHBL0J6ouvRFgyMS4Od+qB1rooKRyUdGTzqRCdn7Q
nhzXO/RuS53TGZg+9UBsO9mT0OaZqpF8+U1l71mP9Q/H7kcMs82LWJ+/zNurfD4oaZqP+4b+lF52
2XP6FCkZ5MnY4GV/4vQyUaYGYZoj/RZeWagGQATt8hvgq82nCIrif53hqwWVD/5gsNIeZc0CTd1H
SJiIzq8pV4JYtJzJeySo1j5iQvwLXfpyZETaT/6MOMYk/o49wWyZDTpl5GuKLPdjpXZZ7HsvHvtX
WlMKep0Gpue+P+jYI3dTDJ0a2NpHeGJo9w/GTeyqPrBl4FwlJprI4w/+9NZzYtRLjdWNHeEydstD
8BOMUjo8WNjcVh35xMlnbQ3QycTk8+shI9xpkZjRm6UE9fopYjjdjqKH0C4eHM7nDsvVB0I0h5gt
ZSypZG4hcbGwdoVBONYD9Up2CJQGiAnW4kKDCfc9JpSLfiE6DR5NSgqVEF0y6EEPDxqyVSg30vbN
bdCZ/SdAq3l9mHissYt8BOPys7dnDGNT2dVLwudTrkxamXmF5AtBwMz0bueSADU5jHoO752xmYDy
oC0LydviegwDhPe1a80NqXCPeASWxTskfgS8GpKtmOF6OxwPugqOHxSgvnnTh8LLTZD3YqasDITj
jkZ8dmKL23FtmuVvANcKWsmH8zYPfk2/vwaicA/xLMjfKL0pYo/ZWXfPSOgHhe3QJhqYXLwSrRFG
4WZ/JSWc8/awI6kHJKajcOsw9czyAGTWsNb0tZFwU+QArXIAXUd1kVf0b+E9P5J4iM/9k52vJAd8
bpNQQrU9IT95XkneiLybc2X+AAQXSJv/Zz2R1+exG1FqQ9ladcsO+E90xNHhpBE0la+xjHPadvjR
HEwvjUG8vm+gCuVHDwsDtDuzAE9AHhmixmOqtps9j/QzNHR6z7GmAVxBG8Acv4nqFk6tY/0Hq0Jv
gjcX6Oy8kkb7ekDBTL7kYQYBMSIizuG/q379vb1RD4089Awa44sHPk/vd2T/NJMpN0fmLg9rlajK
cBfI3d8S5iDy86WplM1t1sx6O6KWBzWUKlESN1z+ox13sWXughYhobeHhFh7pnCJMGubDNCx0yBs
DJu9NnnKkZr3wBZtODR5mS8A/x3XCR2BNzbU9FoCSWbT9BFNyk/vix4Inae3uGpm/yC0lOTHntqi
SJaevVZeZhQ8OZuYFWqFcO7iSlDvKvyVN/AJ2vS1/K2hNwkY5fgpb7gnCc/6bu0XcnftwNtubjlN
Vn0z2jBK+s1qsu3FvCAZdaTwboUrx3Sm+jUw1dnSUXLIZLfcmn4kMukXJvDAhgq4cyT4zWbuJYxP
l/TzsV0a+6HkZjMarx8llZ3ryMjzaQIy4I32399/pwzJAhlVjIBLsGq/wQu/Vz89XGhY8c4FrtNz
s8VCuvxISo9ptMJW+eo3EB910wTN+1xTqayXPrvOwD9FQtoBVMkf7EzIoahn3Sx4F0yA6aEsYoFS
JNLqAn/ELHXFTViFUqnATxR1JBoAYclcETb4993tqaI9330rNvw3WC5/TIBn9dak32QMbtoWGrW5
iXbf8i7Ooyr59Ro7/uD2uIrD5s/+QujZsHxGEy91PYfAGYeXGj6R9Ji7FjlefJcEkd8n4zBTmMu1
7XTyPSgktwbbzSxCFv2sFq7PGKGDjZvUuH1WhGg2JH5bfaFiPd+aWwk/WCddWsxdh//nhjmrgACx
OBgBFYD9jCtYg3bTPyOAxwl1ymJiKIDvS6aLLjAee30HZExsPUMp4foVMv/uRcTb12UoHMDuC5g8
tmDQJ6o6CUEQMMTDvth+I9sjpiFb77/p/DX+KX7xoJ27D9cV1H1pAuTmv9pZKQC45TpJ7KbiYm3W
eqKD4dNvqqjhDBBn6sz1tLomuZd5vbdk4RC1Q0Eh7dtC8fSd1ondaDB1cvUFtoXzMKpMVrhaL8cf
S2jFVoQ0YASMwd7Vt0npjqTO5GaWz1wM4cbyYAfDGpQuQck28NcTS7lNm+q5Bt3ugaU4VSzMnh4x
8dgzfWCJEaC8SQLmrdlgsPM6u9nF7J3O8eYdxMWmxydQJIhH2uZsMqz0zZ6O4zT45BwBu+1pamY8
xdBFGg+wiaBBPCEgQ+/iSm7XfHOA/FG02lROv0iw23D63fFLob2jNizKBr90lz28PuU7Kg86Lxdo
IXMmF3PEO2NxuIM60xRlgeJGMMzvn+K3tavBTihwcN1QZLmvQsfJW1Ejw6m2PWI2N2gZcXUBS+Au
dDD9ubqs/ckw6oGwjY0N4T+dzc56V7ZDRqOcmb5umlXa0Vd8k6SmOCfFUVWDupryDaPUIdqzEypg
4orlDlDrYFyeF2ZM91oJIJd1SsDUcbVhObDpAiiLnmN+4z1v00HX2g1gAJEvRH2LHmryVowfBXXf
HDBY5rtsYyVUj8tTca35MnOUzZqW/yeIgol7C2FFuwbLrvcISvuzsLuOmNTFf118Dab56pjAwHnL
lmBUSvuGa597/aUamyr6A28EB0u/D8m+NgfDaEeC6fKY7BEklrMYFkaceMW0gZH1kp9a08Sty5E7
CfjIv8V4UpkuqnzkZKz2OOXvDu2tbJor1go49WeotGs5WMe93dL4flJ7yZCUz/NSk84S7MR6iJjU
G9S2weUHyfo/WOr3N5QGMLy0bpSh84vfI8DDlWyX9FvEqXVP5XlhjGEGlKI4cQBBP2k+Xt2m1cvh
KBIfkKv82XVzuHKjaBZmkSyhj7J2B7X86wepf5XDG+KhO0p/METsOT2f0i3iD5NFv3So+KPDv1wP
ak0YxwFDCQpLzlSFgMGYIIDueRJJk3gqbQo6bc7Z75hLZdwkbEfLWvxgApXGQjayZzjqatOBl0Xo
TrXrBtv1XctYNh7emTUtnLJeOrAFBEGoaqaUZhcf5E8INKvipedDp1E8PbiSxfEebzbgV4Cs4uCc
1aorjzGJyVvkAXKiKkzQ4AXo1baXvOCF0ljfxv1wbz3E+kPphl0S+L8iRPpxtz1VRRRGLpCTKgNQ
IKa2ODF7osZ+Z1CmIUE8gYkZVYb1wPP5uCA5bnfsEheiD+js03P4QZwdPEiKpFYO+I9xzCeH3EMM
rgT9We0ob3T0KyUaxuQFYWLPcVdOnvtr3P5BcCqHYNKsAUF+GXO4Mc66fUneyXhovaxvdd7dIJVh
xlya5L2jnvz5fSDw5rfEaGQKBRe2vnaK2wIGYeeDsjMgD0myHtNsGx6DMlrEko/2AIirr9ea4CPY
N+rKMkwOGtDzNN7DFayja/3BEaVrYBPp26aVuAuvPDCvikEvok7fMUfL0U/uETPGC0UcJOmZyHCC
VsBz1QifBFkvYCt8wLALL5ZsGCgQCgalCSZ/JvX40IlgJzPkPNa0N9SEsjP7ZgsJR2iR+IUl2ZQ7
rLYs7Y+gTPcMebTDYP3QdVXRMOgiS62nSXcjUzD1CtW3wRAIW9Y6xLKYbJ/pjj6gA0gRMVypJbIX
3fI6AbrRQEMD0dvsAkGP8o5MhxXeQKN2r3l4yKmsHLx7SLlaNlW+/zhuitHs9pzt8EX5p75jiWng
gP2qpTxkkw5BuR5GruC/Rj7WGH9klVR8mg7cBY1VHCn0XlddMk777K2rnNFXrRKN6pbDcEnDUL0/
8rN9XDPA1eWZUko015NQmwpVxjiKjo5IGZkL/VqSvhXuWRf84GssgF2q8reaG6v/q6GJzepGL1ZY
9oUSI0hEFWeKqUhZrhNBzNQxAuVlttTusc70fLriNUtRz1xCmizluTXZ+i/vtAUnxFQErvm76j08
wFpYe2o/y4+OQ2ZqpK+j1c6uW7CwtySqoxzNVrcHc0/gxfFJY26NLfuDOvnKRz6LrPacYUohwnh1
BKpLAjKZN/2TpDoqI+v6JYs1nxjkd+zCq3xd+y9l6l58NIyV4VSKQ5QkhTQljhtJYDMs2UdnTLVW
HIOVSaiqRudJ5NHj8MXQ8x/Zg9qakAEPclzUWJflHkK+9570nIJJ09NcWuzC/8Ru+tJg8/AQKMco
npTwFy57hXmoIX9HaNqeS18FyACJSxOcFl94ADKy4CaftjI9/HtqADtuLNJv4Uk/OTBY/uF4kHq8
rsK4tfq9p22TEr9YSp7OrWc4axwc8y/9VtXfN4/vEnrR7MIi8u68//NHWLML2aXM8v6CWXc7zikj
oE30TQrCDA0LF+v+b4l288XJg8pZFB782i0/OcOUUflp0JUWx0ymajlKTfXh0FkE3jc7XBHEisF3
AMZlIvRh+kvz2CDe0CA1oCW+7LaRgVgZ7f57z2N7irQTJV3dyhhBH+V2vkaLtbXZYkv0I/+Mqgn8
wU5mhrYyxZ+Y6Ve8DCEmCTTDRRU51BzJaDejgTl0DGvg8NbMNcdoa6Lr9XDDkrCJZvERE8qJYE/U
paMRrLog1Vl8Emlj1/qI3+eQxwgGdVBYyLtZWvqSx2hLOzKIU0zP28lXTTRGjcvj3LAZpdBapzku
nssfpHW4IfBeEtnaNGjquf3zHIKdfIFhX6tvVJNG7HCjnwPnkrNfFYBJs3KZOEpgtUeXy7qpfrCA
8FX9s6TG340hLwCc5GHafRAEaJZaF0o251denftZDxqZtelQPdt9bG9wrBqD3oiD12uHMJOlYfVD
PXX+Gx8YBS422QwbpHlH0c9q2bDOS4hZQScS1ui13P3h0Xo9LBfC1plyyb7uN+O7ayBurDvihNOX
TZZLF4WRUnLLY5Oa273vXo7l8ZdctNLAysHlyK22559zitviNwhomHyRo7S4etMfT2q2alGqv2TZ
IeCjFHUOhBvXfbTr1tS10PzK1dt9phtu7M+OyPT5BK9QJE1CcRePuRN68Y9BxDScPiGz3n9j/7rI
4XinsmDxVs9gWMuxGYBVKkxWdFp65ENvQ2yktzL5/sS1dF0VSf+0SdKDt9xjeYdkIfQDiqUHuugK
xYrKSKf9Hex+h/iuYyP7diZ2B3z4AKeop0UGhaN8SgtSmy2uO73HidcpTYqC7xu3WTxKCfy/BpRd
OQfZVAG5M/grhTxClTzcYYaQklN5bsWzYZxDpsZIjZpbAZYpy61Vw9OS+6q/ZSSUxttEM00Cldmn
67YnNoH23YIox/SURo2Vqsnkzfzt8mbml47nBni/pOeotv6SG4md+tDvyiYfnkEPqDFLEnVE0v25
nwz7mQ/fbYJrYvldZ3xbwMU1Vg+C0j9T/lLHT7Sb5Gggx5zOYg/PvrfW9hQFj2fsjtbwZnM825OE
JpNAf04PguBzt+fteebEw53ESlMl103LzLhrziKjQjO7M2bI2FW/J6S2p0V3ZOUqzFKhO0pEWoLN
TeDt/yIqG3oN+LPPDufhK/VuMt0X1dPYxYKKmn0cIDUghv1EidzjjBLkrafsXyCNe6e3VFpE2O5b
5pq92hbJHyLhUiR3EarXszoc/6yw1lH5r/dlLkBO4PIQrwL72s4C3bXEumwuquEtIX7ydwH0xsx5
vx4VWkEEw3kh/JiP78mcWHRazF5r3Nd/hpj5KH4XSZ5MF6eawq1+lc/cqZaHkeG71ktA3oN7F3bn
LgWNOez4hnx6t4LYyVgT8lqzj/P1YYQq23O8RegV+o59XY3wBFx9RqsTNkbP8AOaS9O+xorTCiid
xyDUxKN3Ft/n4gRas3x9lC4mA+pCeSdqu0rElHgbPxzAonmfYKmK5bCABZrzT63wFo8VLDahqQDZ
BgSsZOvWsrexqbXFta6jbuu7fK62ziUAk4qYR839nDXtEOtfF0rR5Ua64fniLAIrlmoEwKXal8nY
jedK1o3EmwyU07JEKpeIWAqtQvVMQJpADnRH3snHDQ1YIJbFVUSWWzl0EcedK9lCG91xQW07VIi2
y5Ya2feLhXVB8FesydiWxsrF1r5RpqNEdlkpphYnem2QU6rTP1vTHEMll0QHNCrRdArT/BNJLKd8
P+NrFpHZlGp/l7U63Yv1lKYfOASCnMfITe21a567GRRbzQEiEWD18lEhJAotXd9CVgkF7emUbXjf
NP+lkl9SAzvgBiTrOrKI849INlpGRhCV51KEEHyn1+J1qb8JUkhDrFV3zi+3B76OEmAjM5iW7Cnf
ejBphM2bRG5CJKWbo0+p6ad3DxSNFmv6+GCfd1O4ijA0M8sL5zyhiIa2BxOBw/hkFU0Z1Gk1mSn9
6vF1nPmnHTNc5RjSyrNqR6CWIyTVY2XLeNm54iUYsvkwYhYC16gIK2oll7t+w89WIszUmNZ5G0Bd
wQ9TsGlnxwHkvgzIWpdE2BkfXjFZnevj5a0t1uNpK+J1n7o68jLAaFTWJ067htdV3QiphKU1RQ5B
Xb+dQnAwAivacN2RAJsCiyzsDXlX/jmaazXP+QKzovQFLvjkHPALipFOaKdzBVQ2e48z8S3qTyYX
Fycndy6yPKMqgVyqWWk0ElD8tYob2ae7Lv/UfcvuEWgVOpicUMz3hM1fd/Nq1099s60gFsybOzvP
c8pvhSI8KZjEqbguO4+nlFqhKUQTS/sQIbpQZfaGQzxL5eYyEEP5EbQ4iChBtDP+sPI337qs9rdO
J14AhtIzZbA7UC47f+kzY463ODqKICi/yezWWLvu5fSlMxRiOesJQ/c7cTc1FXxlh9pCxKq58bC2
h2IUMOKyYBgvGZpyASV4GnU3n2NoHNvIrUR+fpuBrA6F/mFMihcDnrhB9wsHJY5e9gORpjKHRhbg
mRIUyQdhBNLmdxTdIWF+p0FuiS+y80UB+LF43yDV+SAHGHs14tbYruJa1aAJa0dqR6AaAqRYNtbo
lNN4MzoY4+79W6WLUyzSv9wQuj0YpiubtnLSpzPQ+MHRZpH7+jdMU9BZViYMAmOrlk/UVcwrmb+7
qELKWdzDyqRIV6QV2YhsS7mJCiJgYSPCOuphYaqhPg6wUVw/Ze7hkJE/ZkvTyAmbJEpa9RgwXQwH
p5+WmZO/VTbsICUYnz+Venebkom+FcqV1jCbkX2fBCIujJ9JPBLfrJi6GQdR8dDUf0Hq6IwQXFUK
ClDuPBfSxO7NGK0D6hS22hAAZHXMlkgvJIPnR58hYjpxskcEtFKiG58yi1JGBXdj2wAvJ8sFMJ6H
mg1VegsubjQFf6XpMCV4/EtDOAKB2HEodKyizpraSsSWmW1N3HBe42shhSu7sXq/rRZFSxMfU8jD
itYmTUdSk42flbWOcG7kNABrnKdijtoubEvfzDXAIzQfnUvVB7GVft5KXY/ByrihL0U2xKtjmNPJ
8TTjzoIilY1w/yfKXphZjsru1Bcoc6IDgaH29WJ7/iMuc7J8BFj6crCTt6n6+KMv+GZvpOMKcGXh
bpErbqyjfNJfwrCZPGKbSQXahfsHt+xC1YaWg9wzwekBDP9zXRkAQTqTJh0/X7HLJQjQQCMPwFUV
V+UK5op/WreD/l3uTpGEg6sC2EXzmU7s0PZsukFKdTvhgOSxjXOqWkAJEvXsl9BXLHg4u/zT0KGD
u6GpCK+SmKldyN8TIa/e68DWWgnPCusMtSKNSoLFFDyrLKJcgSKqs75JOJT1mcWgdLr2x0rox+o6
deRGhO5UcQIe1gkyC1AEFQG4pWAiv2Cw7q5f4gI/1b4VGsJqCIWs4VvaHvRrEatVovpmPdkNRWRz
zCZk8P8VUqI6bk5GGYqWdm+rKKNLBiVPAWLb5luu6kU/FuVdVBwJSsfJtah6VRVjFOLWz7LF9RUT
T6NMDdPgArqVjSKt0NbK+G7AzTWKV7OxRo96YSygjQinrQUI3YiSIfYVc0Lx0U4tDqLSMFfkybnB
6L46bhKqYngLM2lT6X7cVmA6MZ0hFpjMxfmpxMwHnDX7YeRfIJA3jiOTEl5Ht5uvQYUmOQ2SRDvc
0FeUn5D/5c3soiOrJuyDYIJhhXfyYqk6bm2eFOYEU/57Vpu7rJpwdl430QAly58oVAMY4s2ZPqCa
hfqu21gHQqbYGPyu5Y4xd0u8s4dS2r+ZAbDBgdBkLfgn9OVTkYVIwd+eDEYkJrW0ul3UTqq4sfO4
KiSx2C8/GiDU0V6H3D87n+m1PyGKILX8B8YVWxdMFJ/Dbie6bKQO4o2Fl/QWePfR0hT/zd4pPkR+
6RtIFN4DLpU9TP2Zx+NA/i6/HkCzI3fk1jojFfgp/Fwe1a6X6BtcBOXpC8SfilZg6w9nFmQc76rI
ugHoGfMtKtUd9iJejB8vru7YPkblxbB+xp2D2MrGLV1/3sCBUgbtUQTeMRRHFs/zf2E+ljXWiYnx
RW1k4lWwhXTqD44F+IJ8EylwK26SZu1ofyNhGn9ka7Y+mFhpibdgirL0ljDc4EmA8bIqjgXuXTkf
m0PQRBE61MgBu/8dKmldmXuq/+sQaVsKAojtNe+CaGMSj9ffDX/8sQRBmdWKLdBonrS/tQaZucf4
wogPjnD2WzcGBj2dSk086GAQrstoaUbhFkuBKZHXOeS00Fm8XrtZODKLQ/SkZ518nFLpw6VnO2/0
ep6Dz+0v+vgDtICnUp+rBdfLblgmXXfIfYjPLa2HAyrxxL07mxt+fXxLjQv50mp6h2gu7AFa0jZk
Hb7/Z69UYwHtwyhhSoPW6PHeyepNWNKy8MGbwd26dbU/TCgnjeOiFwwbmBEUo3vSuVTVoXfmCHk5
jYPZpfuEdW/+QoQkNd5crPqTbaLMSs53gCf9y+5pBu68/U/wp5KLtK4jxhBZsud5MLb6HZQL4sBf
lz26xVBvNxaIdNpInIjHgopVZrpmbvFn7wYcWDhEpqNezp0hKK6uqRLhyl6Ca8Euh9H/LH2pnGVn
gm4tXBi3Cz7QpvQWrh+x0SaC3QUMWdoluB35AsYNXFvi1hBJTCGaYemPkMTYnHAkK2RMi7haF0PF
RXUEDE5Io1jRSeAu0a5lEPLbqXnLRnep+F9UYUpWOVbnfdxbhpneynhdK7JRxSX+2L4gsYwpcxIi
S3xxdznlk579NuXFTtrb1prUWzaRmrInV9/IUEw3AogDQaBeor24v+TeiMVplwpDwHcbXyU8CYNy
qRgYHSZ9tNfgx6Z49u5el5J6ylvY9DiEJIRQEwF28ZfT4GG8POlL4Hf97ZNXaz8iHoA6EMINNmoZ
a16nouN5DdJSG/uGpdvADGTwv2FFahLPWKpYXx6qnoiKPfoKsfyIIfDywcBM0Q/U79tlqpKiOrVY
URPaVWB+NNI4tFnutw1inGoycEy5N9F1b+loPX8k3k38+8OZoB6G6wu8wJl3A7hb5s09C+CpiMWH
G+fq9aBxb98aMpJb1r9srSstBVN7vuJctKqJSLMLhfZZ7+e+ocZIsUFQpc7zFecWlu8D7nCuMldY
7JlObsy0Z1vZpeCAFoFrzTPgNRifwez8HLnyLvTUrRmSHfEqxf0MGWwxcGBXsbGCondOTWmoDNgW
dWiKfp0UZi2kRWQU/NYnlV07aCD6M+hV7jywVyXg+weO/17tMZawrSuGcuIZ0QP0+cHPHF9NeqWt
KQ7c87cGxrt0e9J+lspEWc4t5y6BERn1sXJbR/hk2qN2sNyUvUwqSk/vuqJzNQsTIHmui+9eccDn
/vk2OMFZjixzQwNhWq45wvlmjilN9ug+ZdXwh/pVLcHpsc/Pp7ObN0fWCOmc1Q+8p3/TSNB/zPJD
tVe2fpWXPnTahWH2BIwXjn+dIdZtVE+Z2s3xFQWtLd1ogMDaAV6zhPsHc1uI1PnoiDdDkLU+xenI
Fd7EcOklXu13BmvVnLMneJ+DJrfhScHTO59yV/BsWE6IfWeP1+EDNI8L+I7ElFReBtmWvoGXX593
d1Tj44t9O9jPgOEcd94yqV3cV+RkCWNnmBlHLI1iR1Uv1mb/4xGEP96nEIScwAQx8OtLGqC7AFXc
x9xe8v3uQZ07V21l21HWWSxly5mGQ7j4thjvXKzDD1nrA99y1Of0SRmhD0PtEMxCFd2D5qdgEag7
p8C6986AHYrBx1qXRrtA2fJC1z8/Y/1jzWFNWZ6JZPOsVXe7ngA7DSbR0+8YP2AhFu/EMZfZNpSn
Y0qMw13+lY4gPx4CoBeyqIde1UY1/2taDaGmqN5PAeN7YK3+4E3ybgQ+JxSHAnCwo69S3+69PMpO
S2SFTiXmroCQewe3gqEdKlDNx1eFaRsjcoHi5EWzmuY6hhGoQkDrXHwUjGs7v3RX4b0BfFGfc02B
gFNdBJgxEDE3lbKhLyVlxv2DMk/jshNrig62rJF4KVSpSOzq4mxHzoBYBYFx2jvaBmtoe8yJVdxE
xIc2+xbown8jPOAe65uEacRXUq1rfh7Vltds3ZQk44gqN7fpReluTEJG5EmHP+axm06oVVkOA1Yi
2u9j5ApcLxzbGtdCBin4PwNoVWYeDLMV5PIK9U0cSHl7gL+ye/nMVgEaET017B+Sd1GHr2jgr3wy
MD50Pi/YCRL/zYPUohC0l+fIHFdS3dHRZ5ngxdnzAPfpiYcle1F6Xx4iX9y4o9HTJR0C+mwQUmZw
pGOIW4SxpoBeBTPJbLV4xg+pfLFTPbCKC/h7tGlLQFwhUfgFXeMVUuNSwGRn0en83QEcDLYUoNqX
MBjW+ETsOTTMxTJhf4y+8SmxZ9uPlNHbru2Jk4Alc/lJE6zdHz16ozXwDVzxTO3rAu1bWZcB19wD
NaIG4xGFfwiWxEVu50WSDI8mvGtIi8oVopqfQAeQ75fP3P14OCz5CPyZb5Tf58yRki3YL5G8G6bZ
aCFgeFmF6t2EhuACUyW/iu7JyCv9o1MJZT9M1LeQuAvsHkxZdeeqqjZgkv0iqUrhlgyifN13ETbX
qPH1CzmuN0UvatFLOEWk2xq7kfCXVd7DxsjMUzcgR0bsULm7T9QopG9cBqBzGVcYW1Qq3lyfjRxN
qCt1HuSkA4JQg5reZyWwIbm5Jou43OgsJ2ppDO0Cqvs+Y1oITorCLykuJ+t3p51NL5ecnBSx4ZSA
fPWknOv9DQggTOSRqsZxeQZA6AkOD1GORofKCY8RJt4konUvU5vcl8xcEEgMLp8zLaZzDKEf8gqA
eGdy2TT6Pa2LPuseogMImPNTE+j546/UCLlty8H1rQGOQYi963LyEuH3iB799/n1YyPZ70VBLc2P
hCrCJqsLayAlMzLuwXud+9P6GEMFM9InxAiaEjCHVr3u7dGUel4QAMeuWR5hDi/WVClsqxkL3RIG
dZfWG36y8NwXQGa68JwaGULLwyqzBGhpzuaXH6x8q53aCcHP5w3KChbR40UY3klib+wzSTMJh6FF
yszFOu5496Drity5Pn6IfSS0OT94qQwfDQ9Z4twPaJCKD9dhuDCGUOEayr++rcC1f9SHpU04vrwr
An0mGT2LHJpMUsGxyhAflVPPeVNEQ5GlFXU5UKJJ96fo+9AglCgazp7xoBYCKJbh+YZVLMovACjg
Kdu7wGPIDdsfgVebBjLIjiHFo6OkrM7ZTRY7J+FwyHiNRIh7dmInTo7aGi77ehxyfl4qFZoNQ0Lv
75uTxpswUrWcONAQvXxEbV+N8A4DeTU67F91uFaD9ewimTmkvS6/ln3GtWLFmPyc839KsrdD4o7D
K5dcS+39jMUh0stYTxlfWqc6fmXK/SkHw4Zi9UwjFxOha3OgdAuk36+ptzO0oc+MDprZXOXNKO6R
KsLLTfpDjHOADtK3J9cNYvatmRIVXcf3+daLOSFE2c2m49r+CUYnjApcYF7kLZF+myRtZEUrxBHX
grmLAc1nLK1NMjZIXFhOM08diwrYHVLhdxir9sS3TepjM/qK66WUAat5ifwod1mF1DkjWAnNdUo7
FZn0mpHNe2R7FFKt6yRJxnw0QbAhChrmJYQWL5nzsEHjGpIa1BtgoCKSUjJxW0WWiw4GF/UgBuOo
NFqGR/o4DZVqriN/9bWN04hnyHosSLlnwIUhILP8F2Ds0Zr4uG0Dt+WymCVNZ4mLFpoQ+631Vdta
uC3cfoNWfJXPcZ15b8a43DqSfI9BdZl+bLvXYPH+yt2y1l09ujD9L0gSfbvEz3JAZlpWBToJRE/K
3heFrt3Sgls8yWwV5b/4l378FUpzReOk6EzNgHRa9GNgTxaBCtSLOkxNn0i89LtmqI6q36qGeccj
lZaLovIRspvwkzurVLod1KRT+s7TV/tnQCWHNX5wfHLKawBtT6Hf6CmqmPb0oOHDPNeraee8NMG+
qwTTXtjfg4L0jmiu1V4y3Z44feNrE2GLR1fI5PUVQG97X0Fg72iwz0lHmqIolMYwGmUitp5QGgtM
3qit4XR4PU9mGDrjkMxboWGrz9dnsLOeCInm5cbo1m8M8jzhsfZVSx2/JaQ/Yv3t2fBrd4Z4UpVk
QHTTzufBKgvI2nUinRhpvsO9G7M3P9WgdpWxwKI6cMwHma5imXBDwjKAOT2JRxWLBsRUlI/vlFIR
HkhqH2831Z3filS2Kni80Mq4fciwyWdm6vaXVy2Ia7OqZNVezNTIPruzhEM0l3U2fV10eLpZFW+5
9Aq1SdT3Qp1khh4vIllEkfr1+VoqaAh7vWkKd2tm8tm0bYztE5ylbvwau2GdmFz0tabEf8IoaJwQ
K3NaEIh9Z3hmDKWU2+NJqdZrJk/6iOvzMKgYR9rzam0YnkvhgCmAbAkqqRCRKbNdjS9yBShjS1QY
guKnb7khsoqw+WNdV8vFxYXbsy8T6Kdy700G4ZVhahzh1EFlEwAv4JQfBbTjSVDKaWfT4H1qc4n3
D/g7Y0sAjmOiFTH1rFlWVTJvOJlRWH/jzWfpLrE5F4AKQ7wI+AUubc2hFm19s6C158AY6yQ2h+0y
4/9ELvwsLczdkGj0Z2kg1u56bYot2JCHxIo6+iE9VnV+dlmTfh6Zjn/YJZPlGTXTjq7CQUO41mfg
CP+kyV9IIq3IL0TsvSqtpjzQPWSHNDjKjwkSrgO0gS1oRNj8SFYj+LTYrqRzrLqDB8tGgvka4y9r
b11UAb0TS1QhCmCv2g0jjqOObKpERUtBAqO+H7SlWTcoK9VgPN9nzNDiLtlzsSKSFDbioN9xCfeG
A3X0KTkzryKRcoiHxWXUP3+DGiDjCEG+zYEzXXRYv9Eo6kXrVv9zDaeEphUwZumCpNTGqQhRhOfm
yiWLtYx+Bm+wDcMoY7hP8xDJYngyjN4GRHSzZQ1v91qBrt7Ch9wX7h1fhP2pmaguDfsaNtWnt2Xm
zWLr1Ry31keDSEWStxYrQGGJ7DxEq2n/sPTsV51OYxPeNXfKO92hz3i0ySG5sS7/D2Bp4+P6GR24
mtQTil+2tkcB/wXYi7D0lQpnvk8lTLSI+YVsqr6Swv+YWDCAj1bp8FJ8Kocndq9UueWLV91QQD+7
32Kt48tIMmhBM83h8hT28QrIfsFcCayAVH9F4vANr9EeQsQd0HsWuFren3Gb641ORH+uqXsMSugM
+PEXENvy6p/a9vhkjs7b774Gd1Jy+4CHtNIQYhmWTd7TSkhby4kHvEQnivzDfyRgJtWoX6phV2/D
rPBOevBVTMgE/oQeSHIPibtvs8MSBEKxS2d4XWkwjyHQgR8TqAs1sI7WhJxX8QFTUxiFDfzEau0N
z/u/XNlSLEu+8T5L7GLERTatoLSBLqyXtTm7MH4CkLk13f1vgU8gtdjqP7QnqOAs5w42HzCW7Vg0
9tg6C55AzfmjiIS+iPrbUDjeY2IVg/0dNW9VnPIoxLCcTmkCkzdwZ1whrgvQ6z8i/ph9+gSAOZOx
fW74XUz0PI6kJoQoFUM7opBrXwNX2HCgsP4qcdtx/MTdHqy7LF1z7bMWM8lpPWjD++b75xUij1qf
/bEyZhbK9SbtP5PeRnrrZOLPcgCqTwX4tkDC1s1z/g+guhKVouzCVw24bLuxdEM6UpQgQRt3n+f+
Tt13hib8QxLNeHoPQrsPlxV6+1cv0J8uFYUMOmrKhTw+7VxKsb3iscbVjPjCzfbHCly/v729tITx
jtELZzblnPjhgpmJrhamhrHibQH2iRUdfkmhyuvOvRN1rWZsNXQu3360iJhVjiPf7hqlWO4AjpPf
+pr2mhnTu5+lTvn7pUL96qvh9yq1OhBHm3J9zqB7tSUm8Vm0IIU3brquSI80GoNZOi2eRDZ3BKku
IdasziK85ZpNylIACfo5qRcznLk5/jnOg4S3xMgdJ6KZVpD1zxGTe2uV6l79Su0kqIGCrLmNZVST
mdxFtbmpLiaa12YecT9yZsNX/NtBEFTKPfEyO5s9yw5Y97b1DoUuEuzfgaudUASedcdBxOLQNX6P
4SXokRNAFu9GFfrEtWsE6U1c5zLQBycxGRTTDofCpVcWTdaTX8IaXLyu/lRyGdTDhD/vID6ke3n5
/uZrrRIZigMWf2uhm00Fp9m2C4mgWYPog6/HxdQIe7SheWtcpcNfb/vjGtfZvbGHKCDGpUIBSdx5
SH+hp4NYAox8I4PJNbEqywfCgSvdC4QR15BSCSF1Wh3otkJK4OrSeo5glbNLAv6pacfwKtxbWRxb
9EFQYzaKdbtWUk94uz1tv0bGuu78G077KTPWplTmV9btgdE22puavIs92V2m/Mg9fHY3rDfpFZ/1
15qJhS2/KTX/PokRu+m9/RF8u6gd51dSzp0okcMIfoW+wBSlpmYVbEkJZNlkvtfICAdtXLUIj5vp
G5TjGQay43Dmn/nJ1Xi9yFHfjikuXsEM74fjYuyCBIBp/lNF/cBluizuNpwQBUQxQUFZDVZP3Rpk
9SXEFk8PDni5Dg8VUhe4FJ5a5O/QwwrpP0jCgzFk3jWOHXY9tvq/dtYeQXWNc+cbT5AkmMlMmoCJ
IBn3E4xkAV7NWlbM0m4e34g60vzhlnXGY0fbHIYWr3OdS9FRCJ/fWYWlrRdgALTJo0QyciE4zGWj
U6GrClzEjVB90/jmTB5Ghaq+09tJyDRAD2JmewVLH80/A/RTSgUpVL8zYvV0KiA7XC86xrOMy5OS
M0X8N+t4h3JEXyILt4MJSQ0luUpUN+y/YPtfEvYam2XLzP7qk5BCksTzNupALmnCOmc2zOzGYHJF
KPwkVnVh+YhauVQUNQf7VD8WdxBD1cLcJytdiYgj/s42ni5G9tdppevo8Kmk8ihX66qWsT9mUXOA
dUTcS8eDz18Jc94sUktaSquhh82052pxf9CVfL1p28YXXsAG9XkoApbXes/dLQOkE1DNSUvc8dRp
98u61VOilqFL1K5OGAB25HjdeAAG1Z+hshwXaV1QircNMmCoPGBKtC78sFh41UWWwdr8g8xt39Zy
ULFmdupT5QYjiay4jejAcFrPs57u1n2j6JL7Lz5yYMRUS8fYFN9FWTVIoRWdxXeh4MLO99yGJhCA
uQIhXGnkxRjbTkwImm46ZU0Ch6z7mpXdYnBB5Ym7YvuqVOMuj5I0jsktbPIV4n6wEpBdszjZVz9b
q8ksldPS+wEaql+cTFsMcCUz3BIzGKZcRx8tl1vj83aeDwodKTloqppicgyLdvbon1AGmzgVaxli
Rl8hakvcdN3U31tyawafogPeYgaZHA7a+LJX/kP2TeS5tgLGolk6+y/DczoFUUrq10edTqRONqCA
Yda72S9YasbvyB4pXbLqfrezpl7A80j8++8OhgCJKhehWFZIWkuX4gWyC+UORzJIULbC6jygHeRN
+7/qrJ1lA2mIN1xO4dKZT8wfW6BUcZPqtpYda8nw57W09tG3Kx8HTv46g9mXjNMm99mH9Y30e/YA
YyEinMm6HOv0y0fCPJZidhBv7aaQkIFYscslgY2Ks6mQjgbXm7P2V050jV2/lNVHUmNbZhSipB5o
J7n1dTTIK8cw6ns9HMUingDOHeoKH3S2xzVCdN6rmrL3Hykvt9IdThpaU6PcsPrUtJQGtmr4djWF
Dkvlp4qxTqNXpldRdEOEtBv5QLFxUoTN35qT0QImJ0KbnqvrziMzFb7oAf5E1Gbw/X1Z/2krjMDh
JEivBDnpe23jVENyIB5ZjTX2N0UUtnLTnYRzB9WiW8l9zMqgR2A9+NbvmdVEvLhwv+9wnwcv3nuP
z+N113XLusUSB4rGHYIYL8sCmNqnXJNHd0PuT93DSVcts1fgE7YBgRVeA3MtYdYzsQj8yghQEFPN
1Z9A5019K2hy8+WQtiOxMJ5wXEsuvH9G9fPMDc3cdLzFeUZLS1QX7mZ36Gj7FKvCyvY7BNBbwGNh
IRjikJ3zuT8CZ27waWB50pXAOhgpt34FdrnpUOqBbFhfF73JQ6Hy5lA+zbspal8Act74aSRASbPC
Ybanse0vvq62rvxXdsMbDAx7OTe+Z5nAt22EPMrgzL0JmZN3T9YaGMkt/EjEcSHww3yFNKAAqynu
8H+6avFBT5JixzCqtRuz5B3LKY8sWNTyNtApbweZZD9SdX6hXv86SSNqPiKI1I73Cr4Hq5+KDdc+
anYVs7mmoTaPolT3hCOC7TycThiHMJZDHMwEY9pNPw5Dog8dxlvovU4eO2RRAGhH0k1bvN8vOxEi
FoZUgEVL97IMtSfCjg6w8RXY27s3+lK7T01JRlXVNpSiEBHDS39js+5D2NnOBkxwl0RbVX9cphFG
3gK2tCsevbwpXwAznZ1QAgRrzGaDJrRxPsGFwIMRfvzwrH+GGXGPy2Q0gIH9Da8xX+PLncsPjPFh
DiESiDRgMHYJgSa+GVeKdMka9V+07gqZz4NS3KLCKx3za+R0KtSR+SaUrGGcRSBqn3OJmusOTbIs
GtU9eXw2TvWRlhfkDyreB499igCtaHzkmbPs81tedq6gUw7yQ6OFuBO4Vuyl9ZRTZV3/mV6V2ua8
1Nbjm7XHMZ10sDZkXskAf2KXq8ihjxSWJf/wThYKhZ3l2cTSLOLsVVbjfr9wPW9ppIFQ9kC9PlaU
HIxR0AFuaisf/cObNoGkzZyB+tRaRfv3EB5YGoYAiUZuUAvJkKOGb9ErH0KRfO/SaO/OuniZgzbE
MGW5zy/YS6f1t+ZI+1QCP55IPmSTUeXWSeui+aEv+708QUZAKOdXOUqMThYwtahPb9WD12omzzgE
7p3YS5TWrDyXftQhtwHrjW0jT9cpDfQ+/YauB77eyJh6IZdAQ+ai6yrAhJTChnV1pf49U5Uf4JW+
qsNsVke3NJoHKB9aU5XiVuhpMmTsaFzzL/pTWd/yuJxRBx6wKLPda418PYY/ask1soOX17UlcdbE
3iKGQ92nRfbpllR5jL4T6Mvnmt9WHe7XCsbsQfyl43NC490NxjNwy96Mf3sWfROeHOITrcMsNuVU
D7vvptNlFWQJPgnkSL/uryhEbE6XTukcKgT0CktOO2Hvd5XeSSqEHlJvuKOAbqbVKrfz2qBdv5m9
NoPi/w9pUOSJcZkR3CItIUYTJdFHdzQvobl352oJntbW8Ht6Uj4I2IHg5thed1G19pKlpR0lBuM/
fl576lI9uuYw49wA8ShMyDZ0AOCOL5C95iWLUek1FmC69XI48gLI7lj6cP9hP57MXhy+jscASPtu
tWhPE+N5laJiM/rYoduibAOlbhS2dT8lHVLGjQPFJMamb+fIyGV32TbHorqJIVPfnDjuDhYusuPR
A4uTvTIOW/nSnoSVN0qrpICLJOgZTsBoENYlS8Pv3EVcRnUXA86a2BMOSRVHJr4/Iet2jX9xSaMi
Rxq08EbojPYUPmJn5VvKIqK1YrSUyQOqv0Rt77hTqJbCG59CHpeiAYW3BG8zrbDlyQtzYsJqGLdk
EO5krNW80XCmVjxtIjvvrxV2V5On/DUpiLp0ECymhQoD/ILrhbFezObI/439Uq7/C3aGzrGOl9Pv
WI8ILNcxVSLtaO12NC10OKtN7T7wf2aW7cWtcSEbnxgXWrv3JfTQ+SdwDSo2626unsi4JIazsOyk
/TvQChB83U1q0N5VV+Xsjz1+Sv499vIOc217fMkZ1IajXK7RYR7+m2cX0qTDgMR7mLsocoGGZtDE
EpSOFIm3Ud3hbIi5mmJfooy7DPDOOgFTwlwRB+Jybxb7Gw5P58MYroIKTmTPvCEm4zQnkrkxfUOt
P8WdgmO5qWqyiOtnzl8PInxOTVUZGwNyNidtUy7aPC2lsqSjB7I4sQiEAuZKAPeqjaTEqtXricY+
NMldfAoQrp6U5IrwNn76Nzb6DG1tx5OYIZg5BuxTLxDY2AAod5ZGuS6oUrhGcBS2HFqwtGYgvhq4
+sxsPhpIsNymKOHXZ0DqNhtXeLZfwQRF0oGwu14Ay1ZJAOvQXZlLBnGl+OiPqPt/2PjnYz9aWoDj
D7YgZ7Gv7ZKUOHLXmLOyZ+sAZujWeLL0c1J7HPtDYPZRrczAjuDIMx7KQlE1stMq6nzd3KRXPf1w
pYFBJOoP2U2qP4aZTx1IatjIWorxX1llBMFbucOry+9/JUJ8pVvjOVRhJLxRpiuPXinXrst1p0jO
Pc5u+ppBJINXiAddvGVyr3gHK1UnXKOnXF9Yb3oH/oMcwD/ElIEB0OfpH7dlAvPoK14Y1S0q5dpY
PrcwmlmTrz4estJPiHvjYWVAPcJEOk2NFZ7NASba03OD77MOLirvT8Hmn7/kIPIFUOlJBfBQ6us9
yQWpxZ3/SjSFWxcVBF7bYs3zRU/1X55gZjpHRDDurT6Bh0QbQaaLY22wfpOmFinuXeFMEKdHnK4r
F89P0nsad1zFIADSvSNYYrwRAlr/pip9rZ6pbFu0KffpVKYJTOIMs2GERXXA/ZGfhHT4RlQetDSP
QEGl/gHlUGP22+EW0hxmtzBxayfTGt0ww1si7KDte7uaHjPAnaB47xHlsYaMMaFHpylDjW+/hw2a
5Uese8kYyYHfj5FPlr1ulOYl5jEJOvBJfuaNhrNbCIW5TfdA6iOnt456WufJVhHFemNf0KTDmCNp
Nm1lkJy3iHYdWtlmO5WxZnPnbVDp435uStRw9Zw9BoLcTlNN051mXBv9dwJUA+jxrSmnmd7NrzXj
aUSKxe3oT/EWAXnsIAyJ+fjVaPz6ghlVeudQtPpbL2G/UmXl8iLlYDiGYNh/8mizFyYKE7PS7BdG
NuEuNv8z08aWSLxsAeXTLR9V/3ElQrLrG4iTs/whxVMSbb3+XH6f2mIsNw/2KIf9dP6TCGV9oBhr
m2ZCVa9XQDAaB0gFI/pamOWyvaYgDelCUqMKyxdekWX4TQ4s10Ygzj1FHZwnDZHARkef6Vu2G9w9
InAdqwwM/i72dWJFFH5k4lckZXhHjNeowzzrWwmyMf5TdtwgF6EkBvv21tZiyfsAed/8ZsY2DF/G
V2RegXa2VfUJSRbGW8vE1/KtRazGYs4KmqN+ZORTotljklv1KNGk2d2/aEP+V6a9m3CLHMCo1pai
/BMAhrraFSImn/ZymloCCrFYJOAPcrX7ADVpxb+fZGc35/tj8+0gnZvnghH7A2oUOQzXjQWf43dv
025qB9Hx4CQP3Gb2J3ld90IXIA0L3fp/TUjSqRRPCKrGSqMI0spllBBtrIRwI5Pc//CyyUCAHLAN
bPdK1ZF3zQ9UY3qbfHUkkDZ7A5++BZf2zgDWyrUKEiImPVOD+NPHpLdtHjFmOjaPkMH+AZn6O5uI
Dmh3SQWPzcvIoj1Y3fzvi9F1vr9OfIXRdg4Vz3Ds8Iph7qeaUI6FbTLYNPGkgCuuuC+e0jOJC80Q
SmXsacsA9mUhNE90nMSydG3NpzpgtloToSrzFXhFTKJC7H+P1SOFKxYguakdLH2JPtt1LUunh/GZ
zbcQM256SeBYtE3/3ToksWPErl6XMVMIS/vw8fBLZSImNA7qK2eHkm/yklXbcFL+mqZBPyhrSw9h
g2RGN3f1P8wDvh+31gKEqrxixaQQANgySCpRS2/8bClCMMd7hUrYYRoJ4KbTHz2ZDIaX2QrHEoEc
p72r18AFEA2HrdWkSiuuyOGOiMCgKccJvfLN1cathFG54mQG3eJdbKGteH8dvEKM0FuVNXyI3iRV
qMEywnuwiRy0WJHSDB6VuuOT2LUwTOVM56NWB3qfVGdVvaDMfwbXRUy99vmUMX9tNxLi9QQI95S2
2FgGmMUoiVE5ZvrCQ7ieScsJELRS/yYt67N1PBmlr3pND0CB8P2VH5BvMPTN6rXuxvhzPdxQ1TM+
HXWvlrmtVmQWW8mkFVgyFz6Jn66F5c9YW9NV+wmY8v7Z0TzaOHL3G/2AZFJDEVTWq6t9O7r/TlUf
Xr/VDQ/9Z07o+FsfnGCRhoEkQPonwRAe6pfCRSzbbfGS32JCUdEYcJBP9OIxzaoaFAW7WSXqF2TB
CPksNWk3yC7Fy/qxT/maHheVihnQc4OBHH2uf1JXd8McENQ3vf9jeZtr4c9XqJyyLpozebUP6ArR
doazI6douP0/GuyWL+KG7t2/I46a0Kl9C3aelXPrrsrR/96GKwreXxntp9FbcBgqu4L2u7C7E/N9
b1Nd16Vx19OUHuVZmhHrXeHOcxv16zY3qivV69FVVre6MH6ngAIzkvJ+ElXCUCg8fTWs4O/mNr7L
YiCGf6smjzHA7tTah/nDdtpQO+zUbYscq4RZTYo5jNKFZnKuwylRY3DdmLgioKffu60Zvva2Mf36
zEVCQuFyT8+ex6mwsNyZIM93NCpJ/oV8dRRW3t8oqQCdMpYYV15h+vgXFnnbIpgJcwRZVMIxZ2G2
mh+sM45u5lLzJRu91XnSWDkk+b1+xVvkRddQfCx/335wDJfuc62XXkN/9PWPRJOhSmxf2aqBTeYm
AacWiDJvebCm83Avvv2Ji+J0YxTx/bF7BJdLW9FPP0bNQii7ep3qzqs79ApfjZ07LW4550rEHYJB
+0zxbUNgVUmLECy+bd4y28I1QoYfKDZnRQjxvRu/YOU14TkTKXDp4nGDGD8uAxDTyM51ydlsr+i4
Q7snkYwXtdbrZ3ekTxi/Hl4g/EFbiFKznYmRtyTXmb5YY0/V1yEv/OB9CWJDmk0pOQnYWNkuug3X
c1dg2HEuog4AOoB/8BlyJJLOV9HYlCn9U4Tth0HH6h5ntoxpyNoZqLLOLSwxaUHje9JIeW5n9D4U
Ux+SkkL+XHRrdxzV5mL16D7H9RjCmemwR6wkb4Eb4Jr2AvVkmPMdsd/lJ+l5Yod5kaX13IUk5DHG
VAO6XKT6unMkFK/vrtDmLjl5fECRq/GmXtsC4xpFYdxDC9fSe5g+m11GnIpDmkUFyCa7vmGgsEky
1t906d3i0XgZPRwhZG+uLpgz9rmtoUL+xAzHgGxy6v5olaae5Sg5JCeyEzDMscv4FtEPUdIjriKc
8uAANaXfnIqXzRqpQuOvAvYSfi+TgfHIukgAUnnNQexGQwgXZG/Y5k14+ivm3/c1v5xel9i/Tldu
UNI18Cn0wPtRT/5s3QROYQiHpHrJV5fJ/cVksHx8X89jT8GzT0C/sfgEcb3XTIjkiH4t+5V6mQrW
82/ssEOBt+VTP4AtfoMQG/YBNBjhhIhMeEEFaryN31lZTAgK2NCfA/Il1VfLSXKbxsR6PHyaCdEL
eQKdgHtDAZFw4ukc1VVLtuXmhRYl5ZcskAcZLRgxKh/qAhsN8ga27cq1jsP6lL25BBX3OJYBYOjW
4i2ieCk4VZNmjfDMEM4MzdTVMg2LIhk4WarneaNk72p0RXBai0pGdw7I+9EFM3NzX+RxxOQoq82Q
1Aor7NC+rFNG62TTPKl/tmmUKiOwFMzFmJcIODZAuDVVnel3wQDWK6mvPnwFsHwN5LQWrX4EoBgt
STL+CoC4gWAFyZZem3wVduBXQKNGhtCi+fdQjI8aL5wwQ1p/d6o1M0j3D1KEa2fkmdnWIWyzxmdX
NdUcRbbnj1HJhRCARSdfyIQUBVdOoqbj1HNtlHeGOf2YOWhX7lZSwkAoiiIbU6dXe82BtBsBGKeK
3SaY4mLl81Mv9ZLmdPDdyxmADJaroc8h2W3Q5AVAAAl0ah473KQYJlsdfXGFCPRVz+1yiLWIj7/B
3n5AcyGgCRCW6QcjJl9NHm4oYFk0gUgz5MFejA1ESA8X4MuRMbm5/LIOCfYCej1nVVKB9dIZK6ki
JpKIkP8K95B+4Ot3QfQwUCmftzXJgYn8ORTykHhnuFtN2JKkp+ASmKOVJEqTtOjJXQ/CMX9nbpd1
hbij95cmCrcfJecolIHGtjhsWt+Z2hSm7eWsa7491tEyM+Wisz1j33MhFE0oxJoo4TLaU7UwBVfr
i+XG7pspmwRh4iVCGNaw4oUGZsYVh7qQ3GObacBOcR2ayK1B03MyT6IZO1PNCIHvOt+aJNakCun3
d1ly337CGOFcvUmu3fK0P9e0Bal1tqaPwSpOVXCUnXZpMEm/uKpTqHmLaOJ0rMurkPe9hw5pgj7Z
w2DVLmVIg6cU7GI3a+Ijq0ROY9vqYKUXA3S9BXROvnYToBpJbhF8frePafKCLrpnas2NaooVqLBg
OeDa6jjx2uMFwCIh8Vrly5mmHri7bJaMeloAcoF14sjAtw/ABC7HUP+eLCC6f1CjrbEtM+c9HluH
1Kk20mXCC7wHrxsfAx5ARXV8LQV+/zjIFXl78d6mdcv9T7ebofPPjkAWg5czv9//Rl7OnYY5arnQ
V4a/iAyBJO1oi4laAluddI46GVQcySShUsc10aruH70bJ/BalC/srpt/C8DGynBKVSzkXkgupeE7
TT3x5OOsnVmD3PVdEvJs5hmmc0F4tMMfiKISDqfsPZIi6y7ycUpjIxT1hZaf7aP5KRycGh7BPq5O
FJYEYy1p3wSQWbdltaew4cTXa22Y6qDmYzvQAWxJDtK3f16jNSzlBxxM0tq3k/k/tAOp9zZwpvAA
nBD43STwAGPikw887CljXVeRwG8WxbZE2x8CNLX/qtYyKMn++leJ5VlUuH14wdcMvOst2g3/1+4n
rwZzjdLRVwEavsLgDtrdThKtN/G5ovp/AJzqFqH2PLWp0pXGNLK9zVjo+SdDuialRe2fdiXRHdwq
YqTfbBtpJb3SRXZ8NOrlQN4hL9wbswkzLNnChQGLzVQDBOpMTrotVOD8lfnioVaGkjPTtKWGPVIs
f6hwxg8ZLLiL9TtdylnyNJqSLBwI4kk7pW4LMr1gJ5ewaipXFLZmYXv5oDF7zs/LUHfDZczPo0Kx
Y/rug8/1dt7uYfqyDQmx32aEhMGHEQvLovHEQiYZGGIC7Pl/aGaXCPJCVcLbXrp6w/+TBf3km7xb
KuIpGrrmd2YNhyqslGIzJbZhB9zv3IJQoD4kMtl2t9Bdu1Jy4TH+/E21funADMiBiUyWiltZBjXP
kh7Nz9iku71wbLf3sjtmZKoMyLJW+mgDcrf8X/ks85p6BJE+8B3DJ1CybbvLAo+lggMo4vQSrzjf
7KHgvkYGYVuWbspsnsN4VznZWv5F2OS7dTrFd2ltNewoxKiGu936tIOQjjWflVT79JHRZDz6nlz0
7DKSNBEDOqNj9Nhy5VGTrGCv3tLgcNerpNU9SxVykK/Eqc2HALdb0JXgKpKakbgBUwzM+MAcvCyJ
LNZa5vAWZ0vfFKrTfxFHkaPFUqcAWShoQPGo/C8PXXeL60Fh4lJKwP2a0+Q6IqEwGsCsX/J//O9+
mZUf0OuAcbMQuwXEGf1eQ6Wl+v5W8WwWcvAusWJvFfAC80NiWLztUFnf3GkZvgf8D270NEpiltfN
sEYDKbx66DLQZ/D8UMgAybY1SkgxkbmAUtJjnr0fMxA+FnbQelYFNSjrHK97uY8aLkBsZ0c5EP2p
XFNMJOFPyNVXVVlOjNPUBR0mDZF6uu8j3Xb0xkn1+sCWOMqdgEi2m8d7QVMvSkrAech+4GMJ9ocK
bVDyHIrzf84wpWmGjFNWM93N102jog1TtLIJFITkLT9Zj3YqKikZ7GKxEqaMGWN0KvtJFgpyGagD
G3rHGaoDTx5z5FKEFh+qjwPmMQdob3Y/VfAzeETFPKLEq0VeYom5hkG5Fv3D0wK7+3RSl1mqRgzg
zxH4N6NllG4xqWUW2sZOmACbv4PLCLxMDxsf/vTqvrBeETbY5ElnzuJDq+Q8UCmxs0ecsEp+YkJW
UMJ+Hairu3FYAdpYJ+446NoPPupZvFh3vKQzdnFevg4GnjXAe6msCkOnz6LtUtfJ3DvQRT9HalWK
+6V29x6Un3+sSdAAyldEyMLNDzW6rEfRBaR/hQmjPUd9wMFThfkXubxkPAd7ZkftiWsI1Xs6NmlY
j69hHFKMX7aw4XUgHXcjTCILKpPqiZZDAZA57nQIsmNq3rKjo03CsvEtmuhPsQoeZzM39PQpZs8f
4JY8vAKHW9Cx5tLGgp/NJ5rI0qtzouiEMRzdUqrci/gtjpKNUtGSJrMmCPeaDrlzygYCM3zJ6Euc
7W4gEPyh0lFArrxpxpZMGJHKqSI6iVSZeyJPAx6DvGZW/C4umPUiBpYMo9tN0yq4GFVDdR4VdNoT
oM8uiycMTwoh5uPUi3sul1CvBhBaJrE/nr7N9wPyaOPTVJPRkOBZNLdp1AeF3jh+K0Pe5xYekbCH
GuKy9PifiHiPLeNeIE6/le9mUOg4kWvqr2Z4togmhL3TVV7AaVUHRtatyULocLfkPl9giyE6rVln
n3PzoHxkochlxVpeq6TkY8hVvdjrzrqinCvXLz9P+bzbMOmHzQ0NGuKf95SXc6m2XeRK3LXoPWZs
3Mnc0or6y5RIM4aHMVRkF8bmVjx1fQ6H/0zi/V5/9A4OWwK8kSleCFBzdm3VoG0crK9t8kWdEULD
EEjmskpoVe999kaUbiKxY6qMzRbaF6HSnXBvV5dDa1qpRcQ4XzFY2Z2wDCmBNvRC9QXynEUFNG9V
t0VNrUs1/4C7RJp8ZMBs6rXL5JdXHFMQzSQ50FH1EfMRvS7SPLy5VihbwAaf4NIdhvPipou4PjOx
ZswcQXtENxbhWQEkF+DhvrE+4uK8hSJ2xZ/6U1QXkdMNM5I5JEqgyMEWcItAgjq2SbC6Kbkzvoj/
jB15sZsgiUwscek3jOZF75hacxuClrC/4D8Vc4eiF2C83JO9ttncZg9WDca020hDVigi/u72+15J
FrUNUuZenld/+vWGYUn0XIEJtqpbGu2/NkuAmOj0gbv3KsZQzdb9SdgC3rvNTDxfoYI6KXysYdGK
bMHWhM6o9DdVnz4nB/Mz971Oh7bzM9HE7FYyJE1Vyi2FYDnBooXXNriweCf0YoedCOcVK2gZpXGH
E884OFQqiLB+ZlW0zh1qsoRWmQifK9ecXj5mmiE3WLOQMb8u6Pk1RyiXT2/y+CxqJozoIv7PIT5P
nyY3Li+CE2z/eFiBWXtFVqccUZefTE/2aNGBs3i1kfgHHHTka+UdWTWRru6eSarDVbHaXeJTr4GD
+zQwVp9UhSkZcqTJ+HMsk5uNelr4IoXhUSyrpeKQFZDVcfvI0adRHbxJV3xP7n8G6ENoNdz3rHuL
4HpbQ/1esCpjtCnAyxyNUX5ZwfU0mfeJSllsiarQu/1b2lUP/Ghi7KH23/hW5qq2GqLSkqZ7r9a7
5yE/W48ZjmBsifdmeWt8rLPolJ53As64+KB1d9nBCNFFiT9fmUPuSy4Vam1uBHohtWT5wPDc6tXf
m7Nw+a8j4wBrI6fuLvUPo1ptFArsam8RwXS/qerABHQyVXD02oOC+Rf5MUx+Kzyg4rM+yeiObhRT
h460eY0dLBdd+uwuiMNqZzb8wz14IjNucFFf0CWSo2npbXeMspH7lX+8MZ2rI+h+5s1bKZdtl0YP
Ip6Os7qaVhVGCBg3G63JVq3kophiMmSrMQ8prQ1kpllRCwK+MBqMvEOVsIbgd+Fv7MrHR+5d2oPy
XYg3jYdrN2KRBGZqvvMIswGMUflMnCdfAlU+3KHCS6X/VVN4U7hZvE6Eeug8IOONF/L/lsqjmG+c
3fYD0xYtN+Gw5WF/0RFJnZu1Sm7RCQGt+zKFJWCt5GfC2OG4tHmRPWUfhageDba17aUL6rUsMNyq
o6XFxvkST/w8x8NX/2ckTCLtOuTQsZ4taJ1YerpaVL/mhZen5l+3hgE55o/paMrl7V71lRh0uYud
s+1LpVmaktVcnZ+WCwaDOUFNrn45Imbj/MHl57cL2bfrKyynSdRtsOUGn6t86X0RKmFYB1/7JOAg
5otI/BhVOqcGwfvDmgSuNZkjDv7u3LMnJ90hZ5AOZr0QCGhW4afrxA91cZp92eD1djTECS8RhpGQ
2xbfFQEvWSq2Otz0SkTT8eH5XXT2M1f10Jt5tHWyIltGp6ZyFNWkDirtLJ/k/C0yI7RVEPsN+TnV
lWa+OKR4SYaKJl/k3EJP7++YwS/JRveo5o4GU8Qm+IG6gJoW3SytVwtxIdBvpsVSuVU7ji+4vYOS
gsFYBJlkjcrFOje4l7JfVqInFVzT0VYTQIGluoBYUsJMDuxB0k3GD6RunhIZbrN+CwTctzrKIvs6
cOV9r8HnLH51+9hGBH/KnddWvZx6U1J1pFDPZUXj2G5qpVer3fDs1ggv1/mlNS+XY+POBkoQ8z95
i7SIodc6KAr9QAkYqIaFCtD162ikz7HSxPBbcXPQNut1+L5+IbLZh9p78/96Nev8TvBJ564TwxFB
EBs4TTaZd7psH2s3Qd13M3x4dQ25DqMGBwA/REZLed4JGMSUYjx77FZ+GDasp7D3e+1J8jTXffTT
hVK1gPl5z8STDV+j9rUbcZ+mcbaKtiCEGt4a0ZS9CUueCLxUHkEO/Yt30qbu8SFOWwR+ljTqpEM/
FrFBxgSqEmMzbKQ0IGiuX096ULcGi96mJFUjVAQNn/nPPmqsUnUO7hyo+L2oLYyz5LNJzyLl+NQH
QF+zw29Qa+FJcO4yaFgBdjJEWcZevrLcrR6T6vnZ6eAVN/UTIIPGv4crBcfJfIPWWV1yy5Qqct9j
5D3+zhKBJqrTZSMi3BlY21NwDSp4zyLpu+wdc7qmj48RdnyugBm2dD13Zg2omjPQymDWApUOr2RI
FAUtNNwIXyyRDs5BXJNAFDEjkIqeFQqbqgYx2nhzOZe6ddQsBQUff3QNP5HLwM/qTieFWUfqP2bt
D4a7q7XTB8Jy9uMPZd+fukoqGFcJhvud99R8hlkfgsiCaexDvAW+E7c7xNSbtFK8wSRp9ctBQETp
Z06sGh27uBJPG9khI2ZdiiH9MwDhi71L2Ey7690yoNHoZHTAVOvn0kigx2Pi6LZIykWw4emr8q1h
ZSHzLIKQ9Z0w6+8Jf9VlWGNHw6ng5/l/h060edcCkxg5pF8kXb1oVqZ6nYxIlWiNQsws+8/7Gefn
XzBA0c3ib6PL8jdzTTpjvTgEkKAWQNf3Rf1N+PMeHrCuaKy/SQDEVhNkL4cyME0mKjc4jweRk3/0
vSh15yqu+vRJk44Ea1PtNVpbAYxsXTr5tVCbJBdyieSsnKiiuA54fG0OCdfx7bmMtqs/+Ory0LOR
sDdeTBnwxks7N0gwylcrYgRJhl6uGJysGw2TMri3FWp4jzumFRLyof8u9WXOCtyD0ZM605DMQb5E
f//HiAxB6Giq4bVVTrorxGR+4uUGk7mn91z6YPf9m7fbfLb2sE2SUzx0cj/dOUurjTffeznqmaos
48YsopiMvi4mnRYb/Pks+bZbqTg9J9z1q+X6tQKcTOmDSvAkv3QxZ3DR6nUsIYDOXXU9saDCyc3C
bNCvUAz1oZ3rcJaQanvQJmlO/ZEdBHkBKULhMY/ddoIw39CA5d+vod8AJaT+vBBLtnt7XP+ymJ/Q
ILzS3NM/VtzvPQcTVmXr6QgjO5d4huvxpjDJkvKa0ZgseVStuYjGMXLK95M3pkTfWKNcF3IjlFhc
Dtbis2KA0RyiTbUKqaiVBR+tYDKQAz4FdxK8P6e58yaUUaZlOJ3iAYvsJjjj3T9YBi14lYIZ7g2x
pK4YFqHGAPcPXBhmVm3piaNAWFlqujSt0Buhmcnmidgslhu5Q1VZ7mWxDb5v6S7NsZGKaAl6e2gm
J1EjQQ4Uwbd2UDSCPsc07Ym8bYOE6kEL4yxM/r3JQ8oADJTX9m9O6J3H51gvThJuZilEFqgfGCPv
IMto257JAP3ngEAe61mgiZsqxKoswPC7G53w76n+sL9nxoObyt6nKlqaDkAEuTZyBzKsoPQw9XcU
+2BdWaJ4VckZCVQdefsSRNnARwQJ1SmEaCMEA+jCry7zCduXlAX7fh5BfUMzlRX/3I1Xn6cOsVPu
0i/x6Aaq3AZ/wZ38NhdSqrOVPAqZcgLFsFFxEjgCVSssHJhDqMVvgMJRv/nIdxYw3YRWwycLMQCA
k0XLWF2x6aNPOP7cIm/39UrXlvnCxZMq1+VEaq0enuA7AQj6+bhw+wli2BwmEKA2ipwONgMjjiAv
YwYDQZSl4B/aE29aK+d7NOqKuhkvSyMHc6L/mJ4BclcJ5oKn7Ee4Mb+8A+5RS5VxNySRvB74rsFb
ooeIQmL5Me4/9xnu1Rmd1JDXtm27CDp2PwbJuov3rzfDTitRwBxQ9ALlfY1jcSnImOTsbjfZw+GM
klVMR3cdAcxhBk5oNv5q7tSaY/+zVrzzsE9VmE7Ho7cgPjmR0OtRYgxChSYkn+pWzK9MvU8J7Mdt
BpdCr7nE6itqmvleGj1BotsqdNwY0p4TPXk43KP5Ri31Ffv+yXhgTfxknsQAP03jxxG2uL0q1OL2
F3BZ89eE5/O8FdwnK4R0cstrxDKxAW91FGvH9lCepY7tLL1ChyV1u9VRCL8pVi03u0aQpEqd0lHN
Y5rgq2cTfCmIppGFowH1RWujzGpfaVjHAiN1RK4Ll/OavB2nJ7Xdzmq8WyZ9H34LF1J8n4MQMe8V
peKe77G4/EdNDz1WX+fy3Q2+h1aLRiWHeLZBLu22y1wJvhefXrH8KwAJUDcSwpwkReERRDAXzwEz
Yb0XKz07HVeclN8yx8UJw0WukDBnuaMwRyzizxeGJHaRKfGwLTcOsFH4sSLY6GyPD1TrH08yjUUY
xVLYnWPhfUWMeqlr5Y11GuVCGmCD272H7QophcMk+LLRTl+S+7cA8lHRg+1UsPg+RN1oVUGPGu1f
lx3vaFa6FUe89OhuvuUuFmpBRO0kFuN6pDeW6GUu+8PHC1HZJ3tAcnG4uoJxoXa6FJaehUdnK1u9
P/eoPA7Wsjenmu+uYZMQxK12dv9mT0OXFwvVM5CUWOIyI5eVqSNmcbwJjyuHPuCqTZWZcS48FH+Q
SevkswNeLZ7zbbrDoi9WlznLBvtIw3WDsaF4UM95/DL+NSYtT2GGpJij/Iv6mT8sVoubazu9/XVV
+DXAibus1nzegR96HajXosELTlfWaICnaBN7U8ev1rMKobvioxTYH+yx468P1tEDlLisQOz/mkZk
Mr6vsH8Y5wOP57qL7o81QjhCHPIPDwlls5NuMo/iZEamJi65rQfrEBNd2y/Fv1udXLjz+njj20r+
Jktr+J4XSK0jwz+jW2DPdQlInpqxLzcIJ7RLWH7L1MEhS83Knp5lgCSA893fB7Uu6pskvuyxw0ZU
meTO70CwWM49Aix9Cm0WKjTvE5wKYdy9kJ6Q1gEkrMjuG2eaUUeHp8I0IFinjbZAi4w1VCzS5KJU
STaD0kNjNGp62yygwuQjcFSNoLinDkdCzpDXCGxJ0btQLMQ8cQBtIyChm14BIew9ZHGVW2HX9/6w
eYg+qW00+PaTEPwvcuay15U+wOoiSc8Ukw13/18kIiekkH2HhDoXWTbVFu2B0pwFTJ5U5kVxr805
4YR0R8EsktwLeDTTdGTmomI5AwcpalnN7SsO1MAiEJO9aTsQDCIf0Fufo+00mQG7/NKKN71BYS/N
N1p5NkHDjkMUMUti8qYA0xfmriUm/Xh20Kfn438hUJZQBPZrmWbc6skbf9AwOPBTy83TKw3uSGmM
qqwzp6ok0c0w+g8ERrYFbP/WPpPuRq5S5s0f1gz+PBRWS+D95WlOBgZ+PGLjKLQocwi9TeGS0udo
8szCMPSlRwUy7apjszFXuCP8ofMlHXgh/+07M4W2KSE1ircpfUnCe6KyoJ6ZJC8FagG2HzRscQsd
aqR8syKeKo88RcoZzLerOZ5V4cKWbN7xsPZAlsAnCevwuQBM7UIFu1xFqY+k5C8ehwGJbc5c9Glo
2H7elxIuySrpsjdnvSJvRRKdN6Zn5E5TtT37DlHD4L7gCct/kuhtE1Aonyxtj1ziKzjHjxK51Pyu
iXdkyPjFF+3VHHZeDs5Q93CetzyGQYfKs+t5x5W0eo5qn3mdgC423wv4MAgZKqNtye6tT6LA+jZ1
xIDUJboGOpsDQx+Tg66A/UTONkyK42rdxUvdudqseLegF6BxVO1oGlg+tYWJ4G2fvsZ8uTwxLp7q
oM4x2e26Jc8JfOZ9SxBolwDLG7J77UhwpYtTJNUS727HAFdHx8PwZHN5NPeM3QxC3VpuD/A5o6G4
6QX4leQFyE5RoovYLGcptV/jS8ACyKAKaMOLeH2h//fS7P8LYeflD0AVcHUXslRta+ewtDuQk58t
nMZNlyrxfKqVyUtOhvtsp/xsvZx9fqbwEhWAC9OWhg3vKT+bSq/POMIFGnpjXYLrl6ePpunli6tg
JoO0wDf9///WjmYgoyahHeUwHzXqpFc3TvuFTSEYBeFUWl5KrWLfVGLPzL2gcgu3+7OD1Asodq23
VXEazYq33WctH0WXuhPd9kssAZiYiXHqPFLazBch3V8u263pbGS0/a6GZfZrbAYBSemk58ZdVdoS
MgYISvENj+39hCTarzS6wN28Is51QLc6I41BNXAgg6gyF13ORFhr2o5FVVFxI+Z4fY9kyD9Idc+D
C2pikNyYYuguQ5u8/wlZTq4mSKhxzJn8lPV3ba2rhPcHacRmtKSieKfit9Qo8k+KJIv6Jw5yM+Y3
zDmupScCGlbgItuAfXms27lei7p0jJyZYgjn452ixCpKZgx1Lk/IIuxezMs55mFbfYBHtZPCYNW0
r6AVhR/tNjaJDf3o4t75Wa12Id0t0tchLTogB2a3mte1reNE8ZmcnMeOCkR7UqU4qSs4Vn3Ntd94
S7fOfaI6FnHoumdtM3q1tEKHkjxaYQK5Cr1c2FwImh3FMYTG5nrYrNRkrTR0eWRXFeKQMWN7kTfU
x/eqiekSBj6qVBWCAnHgZWOh+hmr4pKUA6aGd/rtyXp0XTFn8fgQnCOHOUCmenE+m+lzeNqa7pt4
ooYn+h3lMu8pcqZpkJ0XQDgi8PAEHygyXIcyUgUAHQOtpuj6O3SYYBJk3t5f/sLK/7tMCGWXTKT6
vIwdTnodqMKdrQwa56GRKcGWFyafZqdq103Cw90My/6vSd+Y3nTD1Lz9tmReBfan2qp++/PC5/Od
w01hRUHwQpc+izZUXc2v2Q9WmWhSiKEpPBq9oke80HU/Z1Y/YXZ/D2mMcwZmsHs2+eoclzM8aVwc
6hBEf7fs1tmGfyVZW0DSC78dwTiPVj7uCVYt3MdrFnjy6hT2B/+cU3Au4BpkK7pvagkPHt4xz9nM
Z7k2BshtEjf7X6JrqTjHqFXKROKDKiYNipCfT60IQlfExgG9L4ly+XQ4DHnCyYcU6B/z5XC3MI28
IYfiTwXj0XhQwxiNA7Q1g9p/PSY/jzEr4DZuyq+LQdDSjGc5f9ZdbeiY4hF3WUb79srP6QEfL1Zb
XIUNLcWmnMhozAFjXbDovQUnDwOK1MHnkcN/id8XEnfu9CRhLm4rYVBm6y7PmXbaa5RcmI5cBwlP
Vp0nP1yDGi75kyGT2QdgqqTRsIraFi7zpTwZijID9py3RWutej+B5YkIa9kA3N20PdKuLhdRiXHW
RiW8HUcL7CHIs8u/5sgjpSykPm0E66NY7ZFqAOfLupGTyR0wtfoG1bYAT6+e8wIQGK7B5g0by++/
EBmU6Otd2sisnueLpB9zDxvmJ1SMlrjfnXjltQcP5Lbq216IOhiPeg6Rn6Atcl2ANNlAsKJzdRW/
SVZGitMoUjIHtQ+5661GV36gzIpc69sF2S8Hw0Il5aBv57pFYUlyeDc+2pS/6t+aoaiCwOvAuARl
Gg0AZ0tQJ0rvwPp64Q/Yta1+XnZIEfpK4B4QUoBreVyWVtT48JQ6pYo9uCTUiqIhWi/IVW9Wy2U5
M7TlHuTIcbwr/WzJ5GcRvyCiwBC09x4pxzwSstL/xDq+8Ih1ZMnSc7OsRlnyzKLuRVH6AnxmtBpp
6hg0JwIxZYk7H3A9pnZ+PKiSTLFvs+NdxHrfrn9NX5kfGxfFOcEZJ9ak2oleNUvwDWEbiYLtcize
jlZhFIQInO6vmeD/ZtCm3L9V2QMnbmqfaQnCudjwg6P1/PEvDNBH9hyEVbhZfY+EIoViD8UDSM0c
F4QLH3XTL9O/ZgKhuI5hsE+kSF/Jmg538EpRrGgr3zbXC8FX3QRE6D1nqMSDoLEL9Ps/PJ2kGe6O
BLs1hl5ZDTrbEY5OsQn/C3YKkr8TcWmMnioM8+Bo5hNTSpeBgP/tFTJMw7Q8PdUc0n02ElZBdKjO
95Y4WAam5lzEPyagTpsPSqo6B7JQoABC0u+WVkjKVnMEELUSHNerUSXDf2fISgALN7UDSar930+H
YAY1ywbe0lIPj2n5kE9UPgLCPqWSqXDxj1QfxgHGDjehEf0qSKxrJRka1NscLP3UplKOutde91Bj
6pTKZ+QzM0Ki4XJ9OfEX4+JXjVRLGFNNL4NiefvPyLBPzwP9qjco9L874LEnLv9kr59Kz4alpn3X
7C3PsTJ/lDHXQT774z52HSiUC4jnogCczaE6x+SIdBcVI7DHaH80K2LefUppM6C5h0T10rW92qJa
wlbJ7tKzXAhvqTwBWbwDjXlmTENMwRXSaCBpbfP38MQg5RVikup9xULrEZxT0PLGcFbUDJkTex7b
BoKc1sZ4hezNG/uKlQff4exCkF1JPbjq0uKhwN/pr0yqHTsNQcKyfMZ1oRvj11SBy3LRUOy8Hxav
K9ddpt2je7n9NzEccuWC7c5tdw99ejcEa61dTfr4S+yszmo44cOB/PotMALHfdCucMHdK0D3TCGV
TmTArxDmjm4XY5BJ6KmHe9q+Bl2eAWOro9UQyBQmZhXlm/2/sJp9oPXJv3deluIDFNLNWJm2b48j
89009DSj0Zqe1dCA9r5xTKmEPDL9BPXv5A5n4WZI3U6Gqf6OqIi26mVvqz+JyxODiFXBVVSmA7ce
I/aiH92E7roWZXpb53fiJXUiuNcrH+u8UK/0JcHerANMRYd3kn2UrfIlm2nCw9F3UKwMTt36uWhs
udFKD5LF3cw9rMpyh0GkAHY1Crdyd3xtLPrt1IRnC14K/000/rE7NEJ2ggUzIc4waSKxihHdLx+C
TXuB4scZGiH0axSEv5HHjVk7wJdR+17IVCDxpfECFYSecgj2+YbyudU6CuDFS0v+5upBioQqb/cZ
gPiIfxARgktrZMGz0SdPZXtKCPCM9Ded5NHfUL8hTkwFj690xeOxzZ7sI2PAzCTpgwkqkFxt77kI
Xwva94NZP/mlVkiYk5Q4Zadg62TrvxBv/iquePpEsAiYSaZayKb3tsN8eCF84nvfDD42FHz2/Cil
CnxLv6iJjnN+qposTQFODtD+CW8xai+BPDmcqhWdTeOmLnIG/5RMpxiX4pL0depQ/aRczm1eX39E
9YZE7JSmw+JkaVkq2QUaG9GQmzCNYos1uaIATFm1VErU1fcQRX8ZVXBUl1oLj8KfrO0HJ9XMjfLv
o7aoU3KxaFHegF+b0scgk1fhPvkIQf+zykmBJcCyypVoqDbTv/xguyddx8E5cSxf+vhYWj/ofBbL
UXdjZrrtHCs2WpwkKtfv2nHEiG6fD0mJrIlRyK9mOSRI2PRIsLqurpHN/R7CLbzpV5DMxJeQ4Ff9
BQZ+wxP+gOmy/NCCK2hkyLyqNhH/YOnXqLZfoLT7r+k/bP8HOwqLvxwKdj2IegC7EtXuKakV4K0K
Lom3+TahU7CMObApEt4fuSC2mjd3hil+a+/UJzMNVorktSdyQZVrhEoQf8XoyUSxcg942l65OZ92
b9tdqYfNHgpnGmNtpQNH1e2WBuXBPq4R9P1zkJOusFNDsUfPR/INh7/Q/Dj13PHM8mfcn+vCAhiM
grLOpymHjY3LD3M8GVRSeytcOIJmPxdGpRCV8v01+npp6+QhXlh9/rg2olCCy5Xzr+e0og2y2MgZ
I6pIi/LF6qgQS/gQY/grXOBH/VxsS5tRWzv5BdcvUmXIaKJ9kWgtJhw3crlMaZw8XicdSQjA6giZ
tgmtAznFXIROBD7kkG6Ho2QzztsjOeVvNm+joe0Xr7wByvhghF1uzMAkSOPyCZ2OceYL/pjr6i9i
BnEnEHYhyohwkHcSBpQodAybOtLhugmJQElqNgcqFgTyt6lKMOqEo8D0UaqWPXIMZsGYPuUOagfK
GEhC5AfzDkqqBKQ4lJcg18GOAOQvS7oJOEub2N5/NA3QV25RNXddGAh2TN/y+VUVIz6jJMyBfD0r
wQSH3eln6pCN8Wez8oPz/Qu9NE88QNTmN0uEX0LVffuMRlRuqNx+Dk5KEdW/vEUgrYdTEgOC8/qF
+F754qyX64fUMbcOCEg4S7dHzPioTX6b9JQk+7iKKfiDV4tw7p7mY8IrOaaVGMXL3u5y2fvR+U7t
ZxsttLPSbk2naaDHC93KI/ZMMCtK1JthaGGrS2Vkc9Kp0ktYQq3B8y1nCxlTuyPr1E3xOc7Pt8+1
G4Gcgf6MN4knCgHM1wCMorg5hdnB3mMwdXZGgqtjYcEyOL6tO+RdTDKQCaGJs9jCLNOKH2YC6jNe
AWi8Lt/qGd9Foo7mzmdrFUvYk90MxIugC0PQkOJgw30owRSSClgFdGGRWIc1lhbyUIyYwAyGs567
Nu+lSSxQObifcmAVwQGmoWZoPZ/MypkqHCa5l4xb9pKpvTNKHseFhqm5ZGuVgPv/Z+pKwjLjhrD5
xO6O2Q/QpVTbse4PAzK9o5YaTNf5jzgl00dr//qXEUMvuksb2iUOOS5u+8vvR5rAZtbCOQjvanMb
2SrzIEv0uI6/aIbL6Ys5x9BfrGfVpvJWC+FsUGdygnI84/Trtn6j9iZe+WttxUH/a3Z0SXcFeilU
NhzYrq5IGAoZv31F8HOwOmf5vbJoUkWsYvChRQPdS6pJ6caEmNvDqrKJh/y2FMUtWkotr//IYotK
Fq0hdRjMdqVnvxoXkBveXmIEP7Ap6o8KE2H0o1CFL8avlso9AfH2u/sdbHkeOZek1TaL8C5wvDLu
4//cwqdt6aZJaf1NF8SZhfSQHBTQpaaaNvivx2B67GjpzyKo9sIzFzWzp8RqsPenvjGLmSSjbFO3
FsMb5gwNamJpCJR5fAthZ9f7XqOBqZys8Nc11GYIoa56irYty57X9g8VaF2YiD43zAHulKQtTezY
vWVB/jbHGanhy8OveXVY+6swVnbM7J3xJNzPUzDu+dDWT+Y0K5DsbYGZMNRe+082VvvMN6DFSfge
L03rItWEd9MRAvwANkYJw545Usuux3Ym5g/y4lnDT8qdMwNTHi38QWnIAfWi+RAlGMv3eph5bR7p
xzemLoZsNZ1rYuCTA5MlRBjdIfRMbjwp89kVJz/1Q+gIBzKer6WWr/QttaiR9uStQRNK3ZDMgpoi
FaS21D+Ztj/y94BG/3xlMawbBr76geqa7axEayjXh6S+nQa65+UKjr8wu96NFSyWw2QLxgFqOKnW
eqmo2zBk5rERIhdgd8q+NKlvQeCK7k+gX4k/OeeclRC5eSNE1mPqA5iHBi5DVWo696jCCe56IRoE
LnnqHzcT8BQ1GYTKzQNcTlQU98mJXUA5WesMtH/OmQLaKsjeDJt0t9X3Ulvxrh6+qRbGxOfnBbJf
f84onEATBQsliZ1hxRZ8F8DuZOnTSTL/vx9OX3nlD/KE9Rjo2YLorVBcD9Q/YwTQrN/KyihTR4P5
Aylz8mbi6bCrVrxw2KVHX7+eCNflJ035UEef7FSoq+q5kRN7iZ5p+IJA3y0NghmbB9B6h7CdT1Fw
ktFF82zoiKtxveShpXchzOvGZqKEefCegrpmE37IWS4rrQXsCb7dFXM8AqgU1YFPe/vrwBTxQe2O
yYmGBv09+A8ExF9950Q8zzY7Cg9rdMEFtYN2qKzGuNtubS8pjHjemj51MxlA1wWKoN+zMv0bk/1E
MBRGBN/v3DvaOR/fnrS3evjzfL0j9y18UjTEsEJQ1I36nforPYwPLQfV1D80tACkPFAexvhGRNL3
/aYOC1UbFHr1KJNxGMuNLVvxyvop+DYWAWW887KJb+OeryCHCFSrirgZCUM/oI9SqOBsY4KTx7Nn
uHiDrSyc6H3cib9dE62+8oHlyn3MSdh5Svl/aC2PMXTN/cmMQHRQ5WmsxwZFBdYXXlQ6d2fqk0Tt
i5eO+QsuZMyFHR4nQ/atZ2+BRGea9M+PrhKrZHpmWmYpGRaci6dknIJKt3KF16BPRBhHgWXUKIrO
ChYimx8GoKd06NzoCRAiqsEdl16b26//c+wjIp9IM5JfyxR3CW/8ywra5fnBneQNiKPsEcfS1ODo
Je1AAmKuBimkcsiXTxWOmgrLFMjU5cX9XbG9KN7+7h+0zGBRWbpeiRQLpb4oufnqjrGgz8Au6mna
OPjeIVqax8jJWP1JTc4T1DjQOdbj0nrhxU/CcEbavTbIZr+ZMygxhvQjcOqXoCZqCi+MlmL2WR9g
Hk9gvnHC9ZjZqXRij7l+GxcQ5ZLtf1xlHlHb4tyklx25J5iZZU1JtnQspASOvPsP6cysWVdTB+zr
UF+KFKB2LXTE7sX7JUxfKtlEhjlyeJXN2y8w0Y2BJM7iPCAtTTEZNxbN1SmcAfIAJsawOfuQt0bD
+2tXjxUBEDZgsuDiU59lfUtAIpT/WmqF1yoaakXrirqTxXULOajk5KhCX944Fvase6/r1PEMjJJQ
9AXoH1Xjc/qaUUsEqd/T+G+zSM92ja49zVVQ7r/l3U6mxJ1A+AH9Hswg/EztGbBr+5CC25N5ZHXA
4FS9ul0RcrETB+e4AWCmawjsuGV/w/68BCKD2GSU4x52rZQWzZFhOoQbPtNK1fjyWteM6FE9Mz5C
GiuK8cQilzDqB0Y8yG/C6Y41BvZu+RI+LHrXhQr5/MBf0qUIPwrCfLUkadFv7gY2Pdu/hulbLVxL
rV33HBGq3v7BLpFcjCmxlutcMK+YBxcx8kaS5yFs7YlAO0a0/KkI3EbIPOR4rjLiTjcCbN5bmNOF
eRytOMGmuwnseNAyhPZgmzcvQhENRkzVuQ07DeH0SMtOyjDj7vxWsOxxVsYp7aHU1P79Z4HeqTR8
sYypShZI76XzPBv6vRbIXxL1C8i5+ED9fLJOpD6MB4liMs3zaKt6+69ffh550rkxdmaqOPemaCbE
jf4gN/A3uANUWyYE1xdUBb/QP7CMTEUoYAGfcEN/lX2gHw3lmmXrD4DjsZ+5MGTwDK6DK8p/WW/i
Q6MF5EqoQxvaRLSR/4CyJCghvCRC5Lh1FqTG6gKix0OA2jEYpKrCM5Sy9mzhjwF2C74RBTfTtA/u
FuVNSpqYPj0I1k1VJme+DS7QfOg4Lvp2m+INjO0ddUU9EB2U4pH0vv39LUorzATF1bDvFNZw8aY2
vMfmm6UQANxzQCDHbaAyN/zfYtLFj6GCTJ6T2ZZlrGMndzv0c5rNVJdSFJ8HeIm4xK0I1X1Sn/0T
VehN/WHgwThTORu9pIcnt/F/bpyAO+ucXuNbC7rU/zEVRCKB/Vypm9topC1bAom0xddDCz9bpKGa
O0b0AGA4WO7kMmzecDNKH09JuZzuwa9D+cJneUZbMA8bG+DqUUVt3xJXp8sEk1AwV5iPBohm0Zgg
xjg3xjYxQirGoChI1SLXmznVHC62IJLSptj96W3fWQB6EBb96vNrF0bWkTgh43v450REd2dfYc7N
IkCjkIH7E8DLq+nPsjqUMOPsjuJX1Z29L0WJi448f2JLcIHtmGnzo2A9O7HFrCF/KuoE2KQHoDXh
qzSsGapXCeCf7UM+mkLB2Bp8JM6XEsO5WHLf+L/Qu/FDspPpu7QUGjCL5wUs7tQYygf8GkMQ+uQx
oen2yePaYV85Z4SnrdNNn8S74c3P6kZDmicb5MpdROnVF5kTOTBS8wxfa0EWcnSrn6C5BOPMnnu+
TANYwDiMMDVabpUjS8GfsWr4yJhgVniQ5vT5HrgBeFERR443nFn3L96GuIytf5DQN7qHJpCMtGN/
9JFuEFlxon2A3AioWTLe5cqEmRV7GqQMplmqEQ8zf6X9zdA9VSVrbV9FZsZfcDzkNF94K/4P4Q8Y
j/rsXPnYu+yX4d2hQqgW2+yX/5oUjfGwoaqMvQ1JminoTm8AU6SzRCs9HFgjsVkCVOkQJcdEKptg
GTlpu+6SpsOEVRo+5B4AUyJWOa9GDZmzFmV8iaVf6u5vgIv2xJgmO5MduVTsxxk7jWAhekRSsNZU
Ue3O39pmpogTH19My7BqkFafvrlYze4W2q3BqwjTkDyqz92ulqHnPNHJVFAoip06yV3mfXpsafLf
Ft49sM3cQxt8NWno8/F6TMNnNS4iCEgEebBUNKGMht5kQYbQPuXC9iSe8wd8XTu5XBsfvYN+VKmL
H1ValB7OvNORzgBR2kXyCDxQMlFLjNLTWC5fbUj6UtDqMisvJf/snu34SJV8CJh8muC/kTWJnp9m
K3L9Uj33g1HuWsCOcfnk+bCnQ307nRksDXHGMORqzp7HwekHjHHNcSxstyVGx7w/V82kCXDJBo80
DR5P46Mo8xO4qnXy9PjjqLf29kpr2N0CfqQO/P7XvoxhPKBw6hoXdWQG0WaEYY7AQI4GN38gDi6C
9+445nGSfW0WQzu/w39ObI79YMldC/vthSNrtmV8+SNGxFH7mgXmoMEsn4EHm+9wPkL3f9VJmNhW
Q7I4Ld3wqiBYEP9G2tSYR6DhWbTg9njZcBrVRiSqG3z0tGGugM390kzW1XEpxyU3K7FLINhPWIzJ
+4AsDbYkI9pocRP3IezTRMgd3Xr/8jIQFzOnpUTP8qapqkuvGklS87ako7rj9XUqIy4ir4j1HxZS
eDKKUq9cNbqX38m81fBTjmwGzC3r/fmVYiDSoT1BtGF4HJjtfTufxMmR8YvG66kolpoXIoQxKbEL
GSOvZ5FPBIW10T366ELvKvnSdzHH2AzyV5QvTCdEa5ZgsQAhmMWWmV8+K/GQtFPw3/hPwJoRALrX
ERr3wD6eiwjglxaV8GoMANjDEOKwVY/5UBdaLwbkV1SqKYQUs5Nl2mEwwekVeHw9BGLt6+nygaZA
5NAT1aUCGk5653EngAK669loIyJu1aNgRBMF9IivrOdtm2sC4aOZ5cMBaUO+kNZb3+hCCvQ4B3J3
NE5fC+OixuQicxAVbImCgzYjDaE6WYusUPLvRwaxCNgYUwn7kyZhHM0cGUep0by9givyQZdZ7/vF
a2c9BYtvx2oM+MJtUhcJ785fWIpK4EoqvJygWjcCp1K9/vpNHu30elc42Zin82nACsr5+w8lQTer
yYZ2CIaG98UgQBXBwyEHnMEzGTkqTREp9GSURjGZTK3/V1EEI/ZmiKWF64F2tiW7x/h5wNf4/y7k
NkPw+/pDBwTK7575BigZXdFOrGxAR+Xj7eowjlCqIhUyIL4/YJADD5jEdPsisk/DUaxc9Jibu8Eo
djNZOqiA8JsiBrusz3KDjSMdqGo3vH73yXcClbTgOvOVAaoStMAuTSP8T+4vkdzZQlnP/iImSU5N
A0Mt+xUsa5BzpfQ06f2z7zhvWVcU2HHrzmkVEhDNIrJlS1fcLPxD68pYufpedwnFk3MO8s68hfN1
C4fNEztLNNGaxooRXm8fpJ/4G3xsl9mFTd7kMkX5KmfVetcSwSAt6TfXamUlwTaYragnH+NYr2bS
p1s3JRuqsYjT3Q287oY6L2GbMxS1ACXbd+knJ0CRpxxYNRNqIlBB8uHPf6HB28RHFfq6694R8rJ2
Yt5o1poL+iWZcqYKyQqZEf8vTo/AKKhvtHd+c+JjPFyqV0bHoTPBKPl/Z0LtZAe5VS2NA8mYeYGk
DUGOZYrp2kbF0hr0Qy9MZ/QyybHzUSnWXgHPs7zZL1kK2fNRJcYPnHQAAb1wWgQKI84xBS0ZyaNf
k0vjFQLsccOCmWoZNRvKWW7RMO1/RuH46sLI4966MprxCiTg0UN483NVbx8Vwk9aId4Tgt8p0uVs
VW1YRpOm5u5rHjOk4580pcOCxPG7bh1DCk14hw4beh6lvX0YrLuhC4lXfqs9gBgivHdvVQeM6ujH
rdOIpZ03+x6xJJRq/cGwA5dk3khK4ihT2Cw9Jtzwgk94wieb5zShIujpeUpclxF2/o9SXHSyRb85
aoJkI30mGAQ9a4x4u9CBI7p1Cvbge2/hbW8DLA0gd95StmyrcSYQ8AeIEAFZ7M4dDE6V4uDuWqUW
QJPgDJfwvwlZ/DBMNkotemAjWEDGNvEipj54HOjwxcznZMKJ+Smd5M6gEE8qoApKk2fwvw9dwgyA
FdSpM6UcM0ifPtSMberwJ4lZRI/2dYl/qELMiQrhzrko80/eSFlKM6jMEfT+tAF3FwD/lFjB+j6i
RJnOllKqiOzl0ONnxSHtfGGjaL86lQIk9wN9AOaGDoPN1KOdrdBdymrH66jkQjnp71ZRu99jDYAw
VGeNJdXXhAyLQd8fV2/gkj3fAG+LRV9LYbSzJGFl6Mva82J7sunLznsViQq9vmic8vMY2FMjES+s
1JdkVC6kWvp646gWl+M4wJ+KojmJPE9J65VM2tYWm2ou14iPiLXtA/uV3NmL5/FqnhX6v/wbPWY/
Z1NNKXHZW0wh3z9AVP7eLGJgguqOzaxQJVygAx7anlKFlkxumQLC6ylqncUbKcdLhqRiiOHuP3T9
k6S2QiItC5J5KmQw3nD8W/tXxO64McMJUtNa0pAHY1AhAvDUZCSj/tRwlvlbNgE2mYHFOovGf/Tf
dRUR8QWWXlGxo7P8zPluUMonZFVIuoMo4LupV8gymzIJ76WxOh8Mlhe1a829c4vdvbrd/hq9a6TB
klgcyTJI3zKR/aIDwsa/mlr/CHpVj8TAumAOuQU14sqTZ8xaMREAsP639fuRC38XMAOkwxBgl8xI
GzwWv9KVDn45z9EGX9O7Z1tV77J0+OuNvl2LOVjfKazNqr06Vr9urrmVGhmBUeWv7Q3zqrQn4Q2B
+6SykG8qRw7j3pYcSMapLlR1UT8tdAfCt+1Drlv2nhF17PJZ1GXb2YUnfGD1oe77aGQ9mkaiYlz9
k5Yvv03voeeHYf0qlwkm0F+EJB10K+md5u22DqqIdRmpkornMRYZ4r1liB/vnoqL/lSH42DoGQaH
bW+GWWvDRhZQHigAwiKIKiz17AxK7t9vc18VQdBGgkd+ROAAPEi0AJnqp3pwQUkZ4tblsuq9I2JX
jcBQ2aekwaoqOHkRU5TV/TMbMdsjYDTxwJ+6jQfkWCUIH0/1Q4VQ7wZKb4u8cV52NGqEuzUaIWFC
K46on48ovHIQWeqYAedWhLeDvp5hNxntr9HPiIUoZdhd9H4xIBhp/Stnj8dPlFj/+Uumv5/t1C4Z
nq9uhOj5bbo8E9X32TqnlHKb5NphSCMhfbOLGC2ULsowNMg1tBhsBI33T6M6nMw+gyuihma4uKJL
fVOlw46ww35PGXJ75ti+hXUpd+yjfpSNAHiFNEg5qE95mlrxwN6nT/svgqdKK/9MYDyt5pTUBThS
Mk7isehQSJJHn9zcMxFrxzKydFaOC67LMVpKolwcRVhjTaH1L8wCd3XX1abO59N8X1sB6TQ381Is
Ym2mnrFLi4fwFvnch2dECs19Bh005GM3PDjonZov4VVES5jjfDeRZDdIppDt2J5QMRE0F5cYT175
HQbT5V5z6fMTKt/LdKVvglE854MFzA4rX20XVTU5eJ+CFpX/UCO4+DOeeYaJWkyQEpVKRIx731Y1
tabLJW79W3154gtPF8XDfSwU2k5R/HaZmFXK2qOByudlGOjkID4YMtKKKWQKQlDhZHqtsFVRNID0
ueSdf731Z0qnIWhZCQ+BoqklvKyDyk+52Rqu5XB+YupNg0bqH3KaXoj0oKxjaAcXlRvjFm9cAmco
7fcVmvaHoSAA50JcEC/frcXngZsFUkDI6JfMObhPU+S9OWrFj0LeaHSH2MleYE9sD2guMbtFjaEG
6WxtNHOYzYfv1YXUta4LZU/beWpXDDePLQ2kcZd0UlehV2BcoH6ofMRQFHqQaq8z681NJfF1a7Wl
do5R676UJ2w68xFFjJA9HsEH9MEE/meOE3cGrwYAfiCI6K9A0ZJAmB2K1MBgBi59roWACPIv67me
iRw/OWIjMP5/+xTFBQThpwvK7jMVA5B3C7RDUWtHh35zJnbq9NvVEOkdY21omJSQkm0rv66hQJPO
ZA4PXVe/IMTFIM8GMdVJJI5XLQrZXGUpgUuC2w8zs/olO4BQqfqxKZEuSt2l7Mz3wm/71EkZqpro
WSj8UuNIwxqQ4DQKF+Irmx5aGE9y1MJBHmTqyJ/Fl1rg0dDXKsJUzh5xwqvqTMgUOiY9i/m7Kx+4
+B+BB0zisRlvhM7++37Fb/3gCsNBZHbkdLmIy2E2UjXCV5cdN92XUrzbUZhAQGFpWw5IlNeHcj0C
2Fa7KwdkTZIDuqBw3rNe+Xv9h8B4Q1cK+oiWElXAFHuEY8AuehJcydZ+Blkm68eP1PTbW86KGJDP
zesXeFAvf7/ETRdPdXVbC7C3my8dp9mptbW7B3UKDzm5HNGvFD+KT+cjw0ePmEI0Fg8Z9vOCQI50
Vdv4erxCoeMfhsGV3th4exdxyQLHxRvgr0PjdaFOT02MZnY4jbcUe8qG+pMve5vUOuT8DhCyKI1U
rMUUy9rCXaZ4yvM2Om77jWuO1/EvlGq2HB1z1XWHnHfN+GF90Rs29qSggMou++77zuj2rH+E+eBa
sBR53naB/UbYh7yVZ21fNebbDkzRVJutLEadD3C8OvyUzrokNsOm+ffONhsEFoWcogd2Ro5s7zsT
RgUE/yM8tSMmvP1PNyjH1Hs8QIsIwuk1lC1vUVXRN2EpJu6lXj4A/9SKzk2FJpHqxYrJBSJYjAgZ
Bqahlkez/QWsFxlb2ebautwjNK87YjT/EAzVyvZ82Go/THhvYUM1Z8i2tSkRnClUU7uZ3muxEC11
B76ZEYaUOjO8Mtcho6CVtX3Kjv/uRveOC3qAcDQhL9KynBBoemajdYQD7RXPDCaa4PHw9Bjht3na
3fGppMjd6ZVdyNU3xvfuFeas9DtfUIQoqmfuR9prbHmd43N9PBJZZ7Yz/Zc3/vNC4UNuHoTD1o87
aKNbRQwwsRbA5rdvYJThhZ6XrQ70fZOljsrtIrwRUqI1XxRl4D/NVe3eGLcuoKDOnusQOW8X5Fvt
UNAv34X/i6wGK4NyMtmcJG5JVHkJM7yJ1mDoA2jM1fJVIzDvIisfHeu/WAbVPwG+bktKAiHSp4KS
z3YfUMXN32bGiYX7CDLfz2n3v+x33YOApWa/w9KGgp6egXfERqfq9vEjUCGvR9a4ypyvCLySatrQ
20Nh3sQs7BCUQWNeEXwTF9e1i1+QwaRvCL41gpiHU5jEr9KTRD553M8lrB0GCkdtFZMpmae5eDEZ
vNP1+e55EPE2Mi630JKml4SGIKpO3iydNQCZhxgV5zais9I/GsME1p485JQhZJ2b49bAn7FIQsgr
OLFk8ZmYvj/QtF2BHD8Arcbo2/1buJIfoOz0oMVd5wVfdSr3KbaOiNdQZI1vS7OnKefWo9Fsvl2z
S66IrZYkaVJvWUyJa2Xcx87cK0sdrm0+HmXbttT1zfPt96vYMoPnI56vaMO90i9HYPj9dvwvYNf6
tZ/hZBuEm1vU/Fzae3LbDu8JXNxjYfmLDR6Wyuy8sYN/qhTDhoItpmUmf2PsOtzhIPsNdonC7nmV
1GbNThn7dsRxonvwqdM4Kx7YRinGwVlDjcK42uwWzLUKgg2c8tHyAFyxx/Sq5ALp7n3MY7Gmpxz7
3LmdsIxD/Q0G+ri7t7JMMNktEWKBSGhDGSWVx2H+cS0Gyknd8hlXSacwtjCjWjAy+vaU5H91Er4z
9Wjk1Wl1SuJrU27YHweIH2bm/sLyRVF6qxi1uuik/ndUiUbvrH4ILNND2VQIrQ6WRlKPUEO+vYeu
WhnSLqVXg8o30XRyouSCMSAA5QEoaXICioe1xmLpWqTgKigt7G09NpKxnC1V19BaN8kFv+xL1TLo
u38KyIFVBvJHU/PEfsgxVDPmYFVTxVXeABC+r9QXq9udIBHz2+vQN3633HQL13TTvGsVouaOSEQd
yJvGtHKHH/Y053F6zBMLqlRfzFSod4RcGtzHtLfPe/AFiByFZM1EL9Vhn1S25Urb3aMWnlPmVjUC
09LVuMwjnC89ExISpiCqFoBZaj0CsYr7vH0nNrs/4fYPfcrGZaS3BWHtrgI3ZX/kY5amvUmzdcZY
h/XwVh//xuQJTTIleX7XXwEzXJqDPVwEMRApZQI+QRXdohmzAjoxuGgoq0YAMgZ0RyPmbwdPPwmP
4mGkJ00lR5e5qgHKZr+aaSRXjvFjaJfpaI5SZ8t2GgnI6uBQCrDGbqHckOzC3LVKNho8skH16aaK
6m95MkhfRAsYILZ2HZAfYBPf4PoQs0oKeh/3Sk/PebKSROQ7bTDA8iDlVVql3nVfPseb/jwVgHLu
fgvKsCeNKC5Yx3Uwi31gGGWJm3l4Zajde3IkWxhJG9v5u1WWjB6wGhY0S+N9j1eh8DFktOfz+fB0
doRX7Fyi2AG1ZNRUfMygq5eUn6vmYpYnUWvZkcMTTi1es+eZpf5dZ2JAjsmwXeoCRtY54taIo0b7
uw40TFgizAbmQzsrbo6MoVMj3jxee08bDzWWy2c0ucqpIDRxaAA6YAAe0j82IrVIxWAQwlvQiIzU
47sI+eYdomqlszZBVc1Gzs1g6OYrD1oiWcpKLfQSJkL7uKSVFg23N1vhHO8XNZkdjcJUN7z1WsAF
mf2LQ+w2spRQvN68qHGNVPHlV1kbiikHX2Zdg1EUGw2RxhdQuFfPIJmrpbLat+TQoEG4Tksoql/B
0Ps3ElfdpRC5QHMYmD6WfxGaL/pJ1So+a3Za2hu035hmbTB6BKbOrRgRQ13gDeaU2nCl53RDb27C
0SMKdUoA+2rRRrd3GhB04yRRE8Uff2ixt2B+F+KSF+DyPARGq9S253qCmuxBm5cAPcEQB6BKtMTM
S9tp+ruZx+TZVUku9ofPHtuzDT0jELtOe27ERGCyjH2Sw0yIEj6QyfJEjDiUX7DrukTEB7jKRpB3
7gNEgBTiZEGBY5rcpR81Kz5DN/T7UJYHRQMnFcsMM4533xulXRDRRVtZPGTstPDWQjmCR1hdmMr7
vY/f6BJsWr4noavYRLYzaFYthQ3ec3TgWo1eXodNM8R8L/Ne8/jXvhUjUT+4W2t5PsONiSSD0rsU
YxDMQiAmxwvQR/t4GlDIfTi59gndREBkIJCu4X+qDg/7NnKKZutyh1Nqi041Gwdnj7FtQOCIS4Mz
mP7gTsqQblbZJcye/GcvDZChAxSqm8yMakyjAkP3xTzbGKxafxJrIVW0PuRLa9oJ8/bzGLXMzWE3
KDVxGIv3WT+VK2SIckWoWeyodfM4KdfTRQXRQ5D0++IkbGP2VKRZzGeNZmQaW3z2R+/86jD1Z4mk
zZwbE32RGE5V+tKyyIKp67Ej7QBtyUSeFAlcsngwn8DTwRTaE5Sig3lFFCqfkkiWVn5dX08qfVtd
DWWeKVBe7lufKfXT1xtDJ+2qtOiZX7FVVd/P3Mn5kMSCXon2uJBWWjLEvlJHwiuwkv+khkRiLsUt
/Ak0WlyV2RKSSGEYKJXmjO/Ory8BlzXwYOIJJIF/M8ZAC5hxzPpBGJmK5EGHJEzcqH43hLSRbC1a
qeH4uUKbYERdJlDFprkAOjsr3+u3SH9fdZLSahCRrVSrMiFevPQh+rx6xCe3VHiMEu/q9hIa0Pfi
NDNWnyhKpzXgjI0DAj5EbzShDnvm+xq124KOSq2WU0q1qwIrtb+TeI5NYEZeKy5GWU7G2sKbobK9
Tj5z6ILHH3M/N82yoYBZnvQw2iVUKGG7YWxw+jmgDUsqyQtMklr04SLxnE+KmiQ4VS9//1adSwXv
cFCjTpciMFc5JLtDNcoZecvExp+XmQBKBqYFXCETAeOhn6R6ViDH6Z8ZUdOo6m82S7w6pNFKH1iO
59gutw5jRHJGhNMG9cGzibC7UK2n212aDnxObQV9k1GB1c6bMZtROAGjcOyU6CI6lJyjlAfPQk7N
5xJejChVyltIEEcAPVWcuF417XaOyq3E+d9q3N60gj06Qbylr4t1pRtN/G7VKpfwB/MjpCbuFn3E
dP6wFPFIk3PNQGaPgvhUnIhU+43R8c2dPCtWHd//3aMT4UAxXjgFW/DWbR1r4cTApkll/pB8d2n6
kGOVvJPpriYLFPXyynoSejB2F2Mye9bmWAjET70AvliVU0rfrPD5y/uEg5bGcMxnsJOR53d9R3sx
rbM/12ATvQHrE8CXltMtAh9ocyIBdXZ3RVI0kHBHFXEBtK2L9sqL85kBd/g+ITAXM7nM/IFW+S4y
r5u5pDXzm4FQmHJNiZTx2hCNH0LXoDB+fuRiDzZraq9VYv/8+SLpwmBn1TeuLudGQ4vhjkdlN6GL
i2K/eNtbike6SZKPqoXMed42D0ZGMlFdQd/su+pgIqTjmoiBTBhh+8ifpjL3r5XBQFF22nvu/3gs
XxjWGO1XTnGk2olOc2tHFEf3ha+1OQBvG0GzcKCkDUjFqpLTBv3mwty37NmXuPCw69P0REsHmR7L
EtftzoqJ5nRaodZRD210wZ41SUgZY9JkczIIaIgj2OXfElFC8DXi5Ji0OW1NrLYYEvVme4jDF61J
GvMHxZwjXR5d2/5euP+hJhXe7chLmTXwakzQd1m8pkDVnA5FSTtwcDf9GHmFlmepHWAYh9LgTLjs
9mq8QQoj0y3Y8LR2qR2qwuWYD6RTnFpRRaIWQTIOcbEECGDw+lQhwNeKRLqMxKF2ywArtmRXYvCi
GliW5ZiAttMzyNC8yC/3hNzc388nbMQV5t+Li0uo+f7UL4cZ3Zll7ylNPcunA3t7+TzI9DFrD6ql
Vm2TqI5Ux+K5EIz5FdX3Fym+Kk9QebZO5MC38yOJNX0zxS2p+BfyIv8yECnfPGy+ldL6V2WWKhJ+
op3M4TyvbtcBTAHIdixaqzLHG0SMTIKZCJ5sKFDekuq+ZkMyU0EGhRi/DZIWCN6YK41Qf1E7+lqr
YCY2fg+6Vt1RHpMFgoAffswcspe3N/ZQmoXfyJpBbX7r6eIteiRPr8bJ2kVqAT7AAMKd3Vq42s27
tS6lKcFjxujkKYCf97XQ7il0fCeyKIJxN9DAAKmSJDCcFXDGHO2J1zU2b8LirD6V+b+8iLNGiAOq
fnzlmx4+uTWdu+gqkIp0/jTRWUxUdIiesDX9STAJtrikEDodnwIYdAlmvIvBfb0GWz2sbWYPXVB/
h9iiwvqTwaLO0wZgwP1LCELNIRQroGrqKUjKjnpC5sLHBdYJ+0mEUoWL/85bjaoQT5oLKv6Qm96n
bXUClTN8K0Bwi7oxtfi6Fo/raXvii2PLDdlWGN7xAY7wcu2Mz1lmE369jVzUSllAk4FZ946XgnBv
PdKR5Li4iBkRfkTINbobCOHBwrqmhph2ERB9G/glVo2Y5xA+yvFO4Zyciyg+r8ZynATKsfu1bgoA
gFSYog77z09OfG47T4cRy0AhJPC+Rsvz9cIAJM2xKZKCZX85WN3wpI9VyVG+5urxiSjRNsBe1U5n
EjY8WaGvpl6Vzdliw+59ayANMH8dE8P8BHl6i7jGJ8foLnJTCji7OFp31ExMJVMwT8N2q/lr6wYJ
cata6aTaKZKc5bR3nw2LUaGBplO7pJ8mWGtN0UqAOdUMpsFdwNMXNwl4ABErPvOUhWCIyJYoODtC
XMwm6v3pwrXmvfnQguUs+FTbGhXqoS+JtZ9HpBViXx8A/ncvLZ8w4zBBi/INH/Jq5xYYUTfnS0K4
E6k3PGEuWSginZVcvkzmknIAS71knbo7eZxN3rz6Vpsbz2NCyyH7Dw/W49yK8nE5Simos8Dy99Xq
ndd2lZdcdJ9G1ZDBCCZicXn2z9sIpiAwrELPXxPTFvtLYX0YtMqpvhSeqGQpEPTTHIkDtKstEYnP
13BhStR+kYVKGEIckLMy4FKlN39gOeYvCVfb6LmCQJdAVj43ySJ0b31GULZUf5aa2TekAwy5iz2v
rkgM4DBwtXKi07E9beMwndnPapi0vjX+5Ayt5z/ohLRq18gWmTPWwfUL/ziCyFX7miC2NOl3uUzB
NQv833hcrDRdTgldPcr1DiPxaOiD/VedGPAWqJ0MeOcHA2zXcx9Kv+CsKsCkGtbAlLwoo/bo+OXx
KPcsW7quvlAAcifmaDaQ+Lwc4cF+YLytBMj/TgROvl3SnsYey6kfkBmX1/AoUx/BvSh7n3vGLkbN
mWl3ZfzkUnWTEaP7chjKV6ls8zaRvyPAa8WBqRBWET2GdLDkhJkU4XYURQHMtHi/pe69QSBm6eqr
eSYVK6hbBEKOkqK7GjxJjftDAIf1mxfMhpEc7ieAXYiWrGe88XzQdTPUDRRh/alrlT8PENQbc7UW
jmPJgfJG8vERph041EijTOs4yk+xahmxj8O04R2YA/PU45US1cyK+JkAPRhP7z2RpUpiZbmTPi3s
UDvHZUZdFltAvUF2tjoON2Pp3IBRkgc+f+sZKxM+lYZH5u1093Y9IlL8O1q/2kpx9yk8RSCM1ZQ/
4UcnjPR5KV7oDawIEJWLwkXswSwkHxl2w85bdfOrF+gnv/yIlxoeBOHsdgPSf+KTI2MpTu/k32xY
MyaWAQ3t0C/LRXTYXZ1FRXHnf/BFS/4s03bP0yNTOn9ay9UBi8TO7aMyIbf1KZ1/N/nLw4cUeKIh
CdWeW3Al5w2OSMYtRAaCz9dJ0Jbp52te6w2wPvaZlJIMXI5Q+I2E1jfvIK/JQzF2Y576NQC9hlnL
+8K3fTGdL8/lpgDnCJh98XJbvFgOzgHxXpE90jT1TfvFOVZCsFW0OTMRecK2M6Scr4nGhFWiCzg/
eU2Wz53klOjotZ7L6wlntLAHk/lFEO0JuG9zq6mXwEAvfAK3iLuvm/y+sNfkIPRwJzSBDJIgx/DU
X6hG+n0oM9UifF+8P9jpKN+f+Dw7QDpbH27/Nqp4mvan3Dlw4PoG0uc5Bjofq1CBfBPx3sUjd0Nc
3FfSQOmpjFnhyUZTZ3rO/Gwu36N3VdH6vCnQUGb3ZPtmsRLPRUZgneROeHBKHMQKmcKcHs8rfBtd
+IgrLjI5nDp7jaKQ3SPGMRzMfStwP4N/argAu4TRteBvKuNxYWEohcyFravT3KlSWD+ND7GzAhuH
QBOHjXFkVlIqnNYk78huxMGqW0/U4rpJ/KSy1Bq3HeErmnaZNFoxQMtZAU/+TtnLYsS9yhP81LEZ
TZflo2xPU0pHPVmiw7WOJ1ANiFn3GnTlA3KzBGHtPiLNIyTUnozXpBRU0jSDcJXo/h8LUmTTfhu0
lLMk+0xrQyVOLk2d++dHZ/1dxfOhZ1hYWKtflIhrbU+t5qcBUfjmpoRQdtyBn3Crqx2h8rXATcZg
wA5/lBhy75FjARBW4bASm7NjI7BG3vgoHxQuWMAUzkU8jhDn6ud5QA/XPvbeHdLUkgmTnxEaDT4C
mG6Zvgl8GHlhWoPUURlfIsxMLdzP+iqTwrIlZAtAZPwwmxwzyliBbuk05SQUtyIgN1LTHncGTyss
NqzpCbsUzLcLido3RQPLzyWIv/0hkL7DSZ0HmQCGxWlKcfAvbAade5BPUaRhF/dQVj7t/zs7WIGV
AkoszS0Jot9jlPhqIKbEbO9etdJC5VaBvUHMk2HejNYnLZKbFTj42Tko2z/kJfDfvtQazEJM/D6o
jbF2F51JMNCvAh3tdoD1VBKPnaCeNAUsUr0a8D6lR1a0z+VCQTI1i6PRoGxjViS9iQlclA9igyJR
30Ia+B8pbAVg0rq+9lPuEafsUthBAF/EmzgTiS/JYqXR9TwzQD6jcms5PaTZjApvi25jvmpfpbNu
tpbYt9zZqFsVpzTA7peJcQI2GyjpAoDpr0AQJTKrt1xA7PsdsGxGC7W/tRNZ9Cy+hHAlTwRWDApt
na0QWVWcmR5FbQEqjFgzkl/nkJL+KXAhG2SYi0xQ0SEwh+XAV9Gmy5+xI+bo2vLLa8EcJV9AkGdA
BjwLWm4PNETgCC8Xfdrp9bnK6v9TWWgdV1YZt0j2e3jcDqQ2IAaxzYmT5ZFcIuY1s8BYy1/+JrHb
BPGC5x/tCoW+8QENPRfSoDy5wg6KqjEEGPQfzV+GsEuzgoweX48TvxIPBWEjRSgYp8O5Y+7W7pfP
+QAvs3+eyWuwhVb5o+JZsw78IcddUwSZQB+NJsmll5EVxINNoUizCteby8U0eNAoUZ2GbzZRzNDh
l6scbiudJ5hcPJe9AaOZRnVN1irLm2Ahxv1phwTB7XSwqFmRDbP9cCLMGmmAT6WeRksNk8JSpy3P
s6O5HjHXfdNgGeKlFRwsfLdIILm63l7frHMrMPMZLNt8PdPjUf/TuetQLS1hH5jkZw3xJWWeyR3c
9Mh2vTRJgMDurXz2JZrmdq80G8OOHBa5TThctsKZn8P9IN48DF8KD7sK3yCLXdIrFrqO6fNTXID2
Wheo6AtA3CExf+iBjJN9mAfinOZiN7wLt1BmZZuOeSYc9WjASi7X5NyCy6Aq6V+TfXxJJgEAxMBg
aimbU4LwtY8IgqYxLfw83IyxRGefreJR3bUMY6/1oBrgs0xJeuc8luAeH6OaB3Iy0RpyMKS4Ir5f
xP0OH8XDgydVhkHQwxE4qC6SUMMqGGM7eGWdKm5hSixCk4vxvhdspKltMgsF3W7M/LdnyIeQLX+H
ZSPcJH5i5+VEB8aLZU5DSq4JjAAHm3Lul/BZ0QncvnD/pEkgDQ3IWNDsC96AhbMhLIooJHVrPIa+
Um6D5wpBREk3RUEwFWQA/amb9ghpKsLGiuxQpjNVW4ePzWqRqUJ9krRVi0Ch/Pj7RSwRQAkAhEVK
1kqzm+9CNQ89eFeVuhN+TSmrhl3EZ3tcM5ybTEandp42Yo7lxNxgVCPrZ2+KKW0ZTqdQigCPjm8V
K7SY7d512gblp059T1Gf3KgMNDuqRr5FbSUPrf+mVO+iFCQlVtQigKYn7dQTYJ8zdgfZj/Kcy+X9
G8gKogdM+7/6RnrgUBG9/0I2EPPf6nRITH/QlAymCCJ4LElS2SgzMttf3NPDH6FYB5sdCKHiyD2M
MSvJpRSSRxlgxrfYYTDKwjzcqdKGfehb7JPSc2PEKZ2WrenNywXEmi+H1e285kh1McN9ansmT0Cd
vccpcORy48toEZao7q7xQKsreaRhxhH0Wom4ORfVS/hmGa15u7PXoyOdIDhBDJwJDZ1mDWQ/ywUF
w3oS3RSxzfiAlR+aavfg+l9SRPR8E9TdEX7Wt15AwNCWH/DqUQeCGHwt1xxaq8zadqwqSVofEIH5
BjEsp8wVSWkWAPofRSI4KHoJNVRCskTXBpkOuxZTjgy0mphXn5Y3gpmf0sY6d9Q0kw2i1jMKsxug
WRy3hcZY8OdMLIMfgDM9gK+yY/HNcBqqbb75Tx5++3yaYH6nzMkwnXCWRNDb7bacMqr/a2BfKzth
k5mcAodYvrlAF0OgzxgX2h7uTi42frCt0rvyhNep8YiVW0uuq8e4hfOcKiAxMZBFQ+NJIbydpcR+
y7pSMKTcRus/xu8eaIi62wmsl1HJZM9XUvElkfkiPQXEvpUCY3Nu7F2MbMmi3yWBzqx4KOUtQq1d
SOdNwmxxZKnHyods6s+7n1AL5GmxC80LCqzkKmUWjWEXm6jWWT+E9BMpo8Le/WK1g8o8PsFOjTqp
Rabszv96lq+bvYSzVEzMRsapXjnpDQjUevi9s5TlCkCE53UUSy/5d65PIqFqQvCDLSkWAdeHvVwr
x6C3NCoWsQxdO48FLkgmkBgcRhlQNpeFApyJoe2vu4agxxzfQU6YzvtHqm57QZ+BZvr84hGEf9iB
XXXWq5rXe4nqCgypP/Ccjoy44q6V+H3YbiUExRxcgP3z/D5p1X8vsbEUcMLyTfW4OiKD5YZPFlfj
GAVh6t4AlXDkINFgwx0g/Ne303xrHM/oy8GLa7RcrCXeCDgPBlV5MjjlhqOlwaVdjry1bgktEkJT
Q79d2RAL8CZgyLgB4BwGXT5yRuCp4Id+nTqughQlS6jNlGz5NRzqeylIvlXdlGCq3hGw8TZXlt+8
PMDDbAFt+ihxm/3TiM/Md8uxsG27Vdl7rOA6SEy4hwfpPf7AfhBQgIpo0dQqDPz8Wo+JBbuL3qua
bHz2yDHjqpT3tqn1PV1RPqkWg7excRNvqQO8OqEsNn/YpFJXeL9FHdGum5VfamOGzd9mmCeCbWbv
7Gl8fczk7ZX00W3Xo7ZGSg5V0hNlFPiJo8BQTVXmWRRzApzumTuTqAZSVOjnkh+Cbg7p7rpPoN1R
tYYh3I2hroYHx+tLugfxWvQFBjFcp0+6JkQU2ecnXT7B6W+UdehLCOHxeLt7GeYwh+mjbGXbMy2h
1MwqVKp5HOodhZmCqG8JeUr2cZkqIVZ3WFxfrLaGlCusA+5zKICcrXQbLZ/xv/PdHAivCeOy1pb3
93FhPlXKaZxUBwqnKB4FjLawBB3WKVQ6dqnI/aHWFdu77RPvXi54KDHAssetIuM18NOu6Jhp/wFm
FB4Y/ZIsCHY/TK22rgjA+ZP+E9HYAl+Qys1lCTIgDOYD5NmyHmAzXfnATjAVMfSti8grNwQYOU6G
j1D3B37edsbBPLBbXWjj9b2gkurhP93ix3T6Y9M9pd6+8TzUtDZBFv+mn8L+w8m5dtv4Ex4BknH4
AT5G/xZp0MaXvmmL/mTX3liLI/PyyUopAaE7jg6KFljfxqKb3nJuJhFAPFbbpjhV2z8VPZ9CwysE
fAQrzziPHIdF3eDdi5E7R1x/ruRfInuU54PwYMbfg3PFD9jvDAaUvbSBeeDlNpGaS5MXK8YbM/9m
vGidVsyAcFtq1dWzGZIeGxTUwwxQUHJEQtQyQSfwtMJATRvuNW9NjMFRFcTweuBi1aSgmAPL5C5U
MoVoXEEsTx2GIOpIRenPDLmKLpdvctLZOFpDyL3AsX8vRUuYDIKCVaXlT9a7EUm4iYlI4OJeiS8h
xoE/Qk2IPbvLPfLYELAsUc2ThpQIRS0yOk20LCjO22s1ByflkF8I1vOUyP1iJ4CN8lPEjrhnmG1w
moxfmohADk5me1FixWFEy2QLlzMCUtfQgSn6UUfGMDFtFpl3veG/1fkZEB6V7Myw6IDxodkwHILT
T/DL5PqDFW5i0l3+RLRQRf5TXnIHuxXKHZfstXfkixIzG4AOqfnL+HjNVnH6hhxkOfSr/Tky0AgM
jXZxzME3fxNxv/aN+ibGlJJ3g0s82ShQTMOwB3fhUgI7p/d7Y+pjGWgYUyASNMKQEFqfOy1nqcbl
vBPO4wPRJJ9GUGb+Av7AnbGt87Cg6Mk3h+aYW7tFin01gv2KxEulBaIRYoTWE9uzlkn9RddW76aO
Zi26TYJUvEkab0M+oiyqtXtliaLOYsf5WYMsbTz7gcN8hdguqlyo7IuBPHXb9HZ0tmqI2hCrjjUU
Fpva/pYvlyuMOfrjCkG5Cm6NM663cwC3bwpuo1JH1HcDb43zgbyReMjhPuv0vgVt/BJgiSNv7Bzk
wD60nkwIFleK9hiGcDd5Xy/dvBGuM3yucvqq12ud2XWfM8u7tiBC71EediWDkLuE4QocGUY7yOjO
Z/9RAh2DGmxkVwQ38LRX1pZAX86x6NxqLRdtWLcq8WAtr7muhV4QPJWRmr3iytuqLFQyoDRBFTIm
mYAfGITBD9tYXhULzNQLs3fEBhiuU6Ys9k5qcOJxmcT0w4bCxEBFrcbY3NloDJGct8+0kCvvYz/0
UHVKcUvboTmdh35r84Eq3Cm8tyYtiLswYFLNbMuPeK6KcrtBnn1ET+s9I9L4HhWbSlwkE+2g9AEZ
PWxu9bJvv33wnchmAoItj+Ky0qX5I7hJBav9wfL+haq7F7q8VzESj3FWF20HtD+Efvvl98GPkvCq
V7IeIL42ufbM7aX+YyyJT0FO4vDFXXuPixKhHX0v95M2ADPJfJLYemYRagr+3+OM//i8XY5jg1dB
80pcRoFFWHR2z2WInzwNWlzaGOR4qpTK+QrSjDpXfRZcw/qr/kIvbHF2MVcVCvmiD3ISO6jlAOVZ
EH6SyxduyNwqvrNG+6wFRrykpZ7N0EtEMDsWOTADceg2R9/4ICMqRwxaSBDj+iEIIBYbHgWB2nCG
67hU/VBw5I/bE/cT7iU1XCpXjHzrq9A+YsC49X+QtBEUwd4BcXl8O3Ev5Qgtx87bylr5kOcuOASd
hoy0MvISKFbvmArW8wJBuDz6ydtFgJKgaXmEqvcoBxRxHNzOmVU3vBA3f32rMqJJme3hAPYw2hfH
2sxva91UOImmSpJuFH3n5/IrlBzooZzqopeDVbPMT00WiTeRJrnUSuYGY0pc4uEfhL8uO70vowON
smuDHLkcJYYSyz5xCCwKwgIgRghF3SqfnAXPm79knkDWSKtbv5TxQeCXU5jTfJZTVuTZbn6CfaAe
RIYpv8ymX35Kw0+rfuxQlSVCbWJXpZrXe7+vs4DROPtOhCFh/NQMg0zT7eWDK4TEi0uGzE7kOgF8
IHq5QbDDUVfcNDvUERs5M4k9h4M3GsJviSshLvQX8qoIltpK6wrBaP+OmWkxF7bxZMzFP2WsBZJo
MJiAfASZ0xPyF+Hs/tCG4wszojNtTTenChvxUboKhX0SBAH6N07nZV1FdpIU6cFy4SdFaHsDHKEA
qL1kyqOLjK89n3R6IpXBO2TAN+lgCnz2F3xRFybZDBKXgs12eiOpJD5oYiqMITorxFsDgvcJkiEn
bZ+kldVtAg4qkrGVwEFTb06g82gvEoOg6V8umvVRWZQj0DI+qnlBf59t9BLvhc1hd/WYdArIbamp
FCovnmDtzdRsQeZjI1kpyuBQq/fBo2vCR5QtguZmw1sf7+9WSX5mapiBIwhwLwku5NSMGGkWTE1K
E13kzhtKEyj/OsFeG+IVF9Jz58YrxC2iR03uZEbUUmtbEtMqE4GqdV3vEXEclBfWu/PzYMLfqTyW
JdssS6a+y6gl3Jew/0Gxyn6MWmYggsf/Ne6rueptYEvo+ZCb0aC8j+xs5VQwUcaUnv1pXO7jm6yn
hsh3imAMSLytBzwJUzlPOPUiYs1/r5PUZnX65Asbj+jd1SwOcNOZIZsQYXYmG0zFJgCg0acLx9Xh
0BGxxfvVAuNXDw+sa6SF3+CvwG2xl8dh40FziyrvKWkJynvLJHjLZUGftxWAKEJWPtqKoidkmLCz
hYakYK4vUCj+270mlllL9Zw5hBQSGfI847aY8QwBBdhS0PRRu1YjZrW34IQDmsGl4ws4r7ZQASrt
ljjJUOBiYnLbK1l9qYG032wPBTmRGdhrpoCw+9EaqDGOYu6PEU2Cz4BCUWhEmt9+ByBFU3kDLR51
2upvHArkq0/q2+kthKrgxl9/VQ58399a1oRdpfDHxoDAh/us2yti1Xz2VjuYe1plJ/LUMfFVj/3f
IilVYCMhZd1u/QAneiIH5Tap9/1reIjzscxCvnngis2fGFXft9Kf5w8aSkr+0a0HyYx2zeLy2UkW
Ov2EU+Q3j42XxaF49F3H+BIw2t9MzMUOxwLWiapy0CMDJw/uYLhq7V+oB2cocH8ONVvysVgesL2m
BkkuQhaxUsnSg4vQaya8K+EsyzmK0Jo+7XXjjIDDwuWHcQ6adMqVRwbVVlK4RoFDMzXZQ/qZxPn8
2RirkRpEX8nRDNg5Xb27b6iBAy+/pisQg+FeFKjoPiSW/K7jLnAjV14dOg54tWw6gIFl5UpCAjGk
1Ssiw9h7rav4yABOZ9HDxM9tBD3wNNo9rysAzt8CJVVH1MKZgViPgn6L7csaskfyVnpyUmMSRfo9
cHVbdmFzmOi4s5yIoL867bWkRDBf1cgn/gLIKOlP0rA27hrvXmrmt96+EMbdV7oSkgxeYPll3ibg
HxQZUfwNbL1GzPamVu3yvbA1S4V5ITROGIf0UcOGxd2KuPGzZiwrBkUOw+P2dPG6RQJKXsh6oXdl
vYRmZOEiC8Ucq2egiJKEoIni4RWw+oFZPmNtagBHF6uCFSSjqREdIsjDylvrnAQb//qH5Vf9bP1T
Sqwq2ETO1G+zwB8BoqyJIwbYBzgE95SxRMeb4d/zQzOpCBHW89nHGGGnIV0DmbPTWC9ZiC9v/Cm/
UahuUDxvjH0hw0BvKDyF52K6WehN1TLcoEZkMDAaU9ewhJp6jMVHDndnFGszgPerebSwTlSc6Yap
fks4yqS0FUtqE9zoSRyiCOuGjW++p8ZEscq0QNBb42BnCey8KFkjWHCBVj0/HtiZK23VxRqIs4Hq
FL+UHym0Snbzngk+02cVVkgE6XZ96X0u07jWyIwYV16RTFLuX33Cygvp4FkjESz8MYMaRF0GOdMO
h6GkzTP882ZNxpoMMp8c7J5ANGKq9XKjw+9EPSplkrzQTEkP1KGXbmJLe1HuDIRCW4SvmOBLZGLI
CNTSGBL6v/lLLnpA1YXwhZLTi+6THPR+W5HgbMEQxukSekox0vAFsXv7kpEopcnBTVkLJcRaLATY
+DH0QU0ntyP7MCjJ8MM6VozjAvnJXeIVWEk4cC3c8D5nlUGEQzF1IsA+9xsYNrfnRUf/lzgE8T+f
6/s49vdgJrSHqQGtom6EZebTiqNh5nDZ8Ikq0lvaZLug8iMWJG7kPMd0bDt+h1TUdcYVcZDY6RzE
5seIuKrRlQx5JZxlWGfjG6aOgKh0hiOBuBFwrnK0JafM19n4RupRbcEfBdF5GTvafTb6VarGL+cy
MNwd/WhtuYzTULTe4EZwbX3xs7+Lb8m2NIBu4oEFPxQilAJVbPN/hMDZ31KfcjvF1WqIJ6nf/MWN
HdJiL5jjZrSRdWWbABgv6Vw2iciw021efgmbuZWjhQdT1WN+Zmm6uMl99yoV92XavUI8qPXVViA0
t3RrYpXWtl+P37+HblTePI9pjOeg4c+/njWJwd6bCaSgogf3RVEGRoqzjBxv0KV/ZRNxzC4PZslu
srLBYBXco/AikELKLRzEHd0OlV0vSJPfnc6WJid/Qdgw8KMVzMJfD7FVq7k/ccWfDPPUh6m065bM
79hZ52/zG5Pb0Re3drnY0ZNf+e9ivBMweztueFHa45WZFYkrqBLu7WzQD7N8kQbfVQzfqfVRfb1L
4NYi8jRgka4A+biCzE06hHyfG8BPmRXVMasdVwf8sgi6eEcmwEifFYln1PpftiChUbbLHKI7NkGz
i1C2Z2641h7LI5eM5pSjZHbiolmwMn5g15WcCdjtJpSIvbOyL8SONWu8Et+R9XBK3eo4ybtQyRbz
tLt0PsEZiuzLQ2ZJSIp0LMS99a7nM1Zsr47fjmfYdWTatKPcddckoHo3hwMOdO6ocIqOeVSXyEE+
i/a8BwECo6fY7G3TPN0zeOsEDX9YluMtBqljP/6Kt+OuWekf6+7w28CGzOPekvnqmHRG83NH+Ps+
WVhW//mN/nwju3AVrTP5CQGVseQaqNVM1i4POO3BcqBuI34Y3lI//peSquf20zOdMmryDZ8cGFSr
wjLCNlXTmWypWacX6OyXrZg4nU90EjNPBIgxUkNiuWLdYApQPPbkBZPnncRP/gPKc+1twIoZGRDB
rTqBTOctgkTLpWCZ3spxcdn/j6x9ExaopEWyi+OzErNkim+iMh+tWQmcR5cvVJr/egUrvfolVAkn
wdk3ZSdtHBxFVFVX32JLCrZnOJoy2DtadoeuxrGdk48bh85PzVacC7xE37uFfGzoD5xAc8ncT5+H
ToVjlh0wqC2uxZtPhxAhnGSpyguvh5l/RWVxirA3ZDf9aDxnEl7Zn2wXulh9IfWUwfy1KOaDBlbz
wAp8OTNQZTcaujY5tlw561zdPZ3TE2W7KSjtRF3rZomQPRoWwhDuGf87Z4dYeSbEkpxRD7o/pDgf
xp03Lb3IEFoYVzM6OhcHXTNE4bZ+1A4wxXIgTNT7MP+oSQYxdxRISfuSP7TWCzxDDluC9FxMmp2f
lcebMcJdTummIsS/3T4TDFypuMQESNeLhxYI8La2xm42wRCOCPmU+xYUDGETGifUWJxphmQxFa4a
s1dbtbB0JWsWotFHnUzL6xCvBHHNEaKVvWZMn8VQAQKHKH9lzySm/Joxf+3BNa7d2b9454cdJ4JY
GxofbJA7KngAWD7ztHJX+MZVLzD7qwFdECO8Xdt7CoBLsIOxcFneeSiKgtkOHCsSBF4zPgo88qN+
xaFn4RkVwO6dqkKpPf5vFyZblmwBf3lwrxoHqUKrl3S3Ya5tJAOYjPYxv/jdb2iM0ZTF6PZaoFXU
1fVNStWtogYgmQL5VwqgZbkcB6SeU0+Cl7kiS1KqZk0yPq2LeNg0I7OckhyGfqcNygEfFvCGOHJa
SNffEr7f5WdFs8K7Srj2AUw77vdI7xYgDuzDMuYMAKvJIsiKuwRw5twXRf8Vf+QxZB1r6KDitww5
Ho1Sh0R1XElrw45wjZOGxLbzB0u361JMLjMdLGW7ilvFJICvni6f/mXkKEx5CIn1Pq3ijtMGZEeE
n6eLeDiJTWISSnYYvFgp4+fs0HRpQqCsgbCb+DzRfkKIp269b+/47dSeeGQnLxNu8bBT7QAzEEkh
P4Av1qQ4kASvqSPRSHFbuLywdIkz/FtMe3p4LW/XTUnEZlLfrPLlMK7p3p+ksiWOQoBPF/oniuGL
t4ZFYSE6lZrNoyw5ZCFV6RHKB3NhyROeDgbrq3gRdTaCCv0JCrSGLhrRT9RstIMMwmC8uELH29eE
8L4+WXd+GgKRbyxiDomdxb0Oj2WbPr037VLlzMkksFcVfWfVYLE32rGwaIf7gdRr/RkcfTwc3Kml
u/Dp1787cvc6P5YUdjGBIb2liTBicWV08o++4DpAEj2STGDTRECwpzJetp9WiDYfQbAA8cdgJqVF
y0INPo9g6a4p2PX+zQt3wePcmcJUBUMTyaySYD1uPuMmU36heeXmU37xNIYEcwffJ4tvfP2e+O5C
Jw9Rj4+JGfg5GiQ7zlAXsu2takeH3/5z4WCIZFeHSCnBb4nXAP8aynn07v6wyYwdUtKduTA23Nl8
l1miB0JMjaPTeYT0gmcxOgt9ff4h6XWbuDPXFuGWyPuUOCCmchsRqOJ+clGiHFT551aVCaWv3lKh
vgp2i24ngXnSRjkUZ+/bFgIMuy6ReebxVReSUEu0B5N7C8Rlc6Yt4JX0PJJ8v2yLzjDPruyMwq8M
OVaH4vaCicL45h58MBOAWiMqXhKAGjGDeggo5EXGBzeX0PIrMRgTZEi7o/biG/Cg2YxYteoWsbyJ
a2mcTXxW/ixmYNuvhSbSywro97Wmf25Qzo1OoJja6l0nDdmHNncQTXn7bgJTNKzQCNgAeUCPZpwp
x8pdseJmuXpXwLTi/WqlCJ2WgFOw8cVqPCMyp6MGYkDrtlDNsoV6xl2LdmN6/JGAju/nvRKAmLlI
l1UEpAuP4e0ZABRMHh39LBfbxuXH2F0Sn+00SL+ZTZGBMus8uRYf43zSN5LZn22P7aIQU0VXRBem
f3OWCBS/Yu3PccJ8+qYhXNYoE+GkeETbV7lGs8+GsxUKJeGxyGZXtLz9iV4HRK+2Ch8MwwLxc/p8
GAK+iT+Nse733DKZ7TSUtwfHZT79uQs/0UC1cZ1rHj5z3kCxlE4o0WEDxAIp5p1RB6ZFUOdho4NI
ti4/RJGs9uOokgVceW66SsL4WTYvK435G6E1V5ZS0lzxsCCapPA/xIp8jfMlpa1iBcrrmVUNNFfn
z1dGKVoP6RRwnkYMjCXm2oXDTwAJ78fMU6l2ctgmyazCfCEMMdi69/uDUmngZRgnhwE/pXTpO9AP
xhsykMNvbFW60QlW3wSn8JTrmxn1gbRFmpZsGA5abEcEUMxnUCcVR6APRbaRfTnRMdBjSV9MUPZC
GwtCbwT9ijh42xMi2hmL4M0DPGkFTES5A9qG7mkfaxYXR6rX+f9X0AY7Rnar6A1Sy9VKtUIFIh+m
X8eA5uawvOP17A0W21vSPfxBwildhTlC4df6bHyrdR0fEW1wjHTTNWYBA1aKDqtE6rXSk7OD7fPB
sVSuCjjTLxaOghiQ+2MogNHpCydEUOhqvvThI1f11OPhSpv2QsOPmtqFms3XayiF8wp+wgQgGxiG
/964/KnX6eAG9le7HLEUf1pu7Fq/epmlZstD/nLMnITOsNl3s3MPYDMSVtdmioz5omaKEq37i0fx
Zg4QG4HxJLvNImdVJ0Ep5UDegv/wyK3D1k15U9ZXiKIm3buv0r9rmqkQcr53aOVBVYSjd5Zn6Obq
sjzzTAik9UcnG/9u+qL0VneaSNqFZjbIcajyJaUBbIg6QEmBe3dklYp570lias+IV71WVfjE3Bwq
7SCNYdWHbYmA5ecWdveEXwnEcZEG5ZcseV4hdTdpsYnFFMHdMl1idFw2CHjAgN5GY2yKMUIqFfxd
DzDA5Re9kQ+La1hE1QKMwxSwnBAHpepTY3ALeUQxnvi0/fcFlfrQdPNccGvRsSnuvSb27z90ODuV
y08lG5nKqrf+1aFALPCGj8axNivcsiSSs3R1IjR2kBjKrA4Am45OPDbP3h31Nht1zIAir5Ml7qh0
3TVda7royUfRNr8pG2RaLqFWsL0RCNxnIeMGoJAe+GGYE34CjqOJYbEghCxEfbs+mtw6U7Qe7VSj
iNiqpKTe3IvMrSINIt3aSKLt/lLv4etgShu9el2v42SDVEE1NJAmxRtlu/S9jE7z0MAJFpGUL+NS
j7P3o8xtRTX2KqIC3imHl8iJewvMfhurCpIEw+ZKBjv03xVuvVNp0EkiXICKmUQ35qrXN1Q9G6lt
jdbFF1+KK+IHK62IkivDxKjzJXHrJJsHmFa9ieTqXTuk5aaa1LXVZi5asrWLmlw3q2Fzun3B+TqT
h+dL8PlxWl7oyFUsjq/jV2ODewQXm98neSjF7efFX4QmPV0Hpk3dBLJf9xjgkH4PSfE6ZdhZbSKI
+o9zZcj0yykI4dVf6mRIrpn36LtpHEYu5uzJrzLSfA18C0+fD5e4i1wUcr5rwaWfqohGVcwUmYC/
C3GPi80KSwzVOhYXKs7gJwDlZN/EMSFqV/594k6Wecu5qYetfm804jjanEDQqTVJLpnMNyChWqZL
e+jI6DBpwtmfMfYNBmofJVJHicy/KsqWn0VSakl6xJ/rP7kdvxlDfJWuifJCRDcgsT/tcJHzY/pa
fwvZ0FKoiUUgPS7Gwpr2IJkivDqHHPaSZ1a2iJ7yL4gmtTSEMhhGR/sXrOw6tLkn5jarLnWs2Fld
S3DXY3mAHCxB/8VxovjwgWrVmKV+Yt/VmOQ6pH3F8jk4Pg/2JpxzJImp3v8op74GcUiTf1KhHfap
loPBqgDoyVUHzT7PeMJbYvN3vpwYhNoa+TFIIHK130CZggA0LQxDylHEIUW+UARg6hdHXAqo8LQo
cNR6/2iBFjM2FJpqFQyO1QcWc9626NWcU8HreaS1IwbNM1bcuaDDWHxM4Tfm1PjspJ6g9NPSRWh5
yW5PMM4+8Qbw6IKxtengGykU5z6JnXLWatZXv7AMZ4Wqa9iQFeDvIspCn+8vszkdZ4NoR76f4A9b
sxIHGw2OVZ+hC1E44FuS9Pay5ycb8neZ6hfDxPp8rb8LsaESA1cxIUn58YlUITaVMt57AwaCgyk+
Kib9oAkXx4wXThW1MPHt5KN92tyP2gv8Fe9KqzuHqiwFmN2ZdzlY4GR6dAbo2fdEQJrcUzXKjJPN
vrJHEFeHOI733ouEE1kBkntC9WF335sHTmJspBA0qlew5yDvcR3FpkPMOfTiHj2r0W6DRjkn+NgZ
cwtNfa0UhTfueyODP2wEFm0nwN86jajoR+Mvv05/Qi7DKhvFtPQ0VjeFYMVHrnPEQI342SSv+1lG
jTHewn6NuaG0jCpPmVq1NzSQrfywQtQhrunXjvWxr/AtES/QZuHy0bMwDtocDy+9cvGyFy3VZx2d
2M6XTGs2eFd7YrZ6T6i/iAOznBnTzoAC4siZIpzKeTM60cSPfHRcA57yc+a4AS2GKDQ0DhvAanQ/
N99KGUQNGAL3XpMpE6kFI/Rzwr9SSeESgWBqk/vOi7pvi4hb8KyVOzRDE3FJCV9UuqKkWL/ChAVT
8DwYCzjZjbC4+8JWRmMk+ss6hw5r1WlNVm9eXFa4Ut7Q0QGDzb5C13Xj1w7U8ik//jkQlOC+tETn
WfS93G/mZkpC+tMqfkV3Zo7CXuY5/K9EhcaS8b+JfNnIR35E1LYpoQuuIqqWURX/cj7Vv8Am1Lwj
I6lMhZq2gJVNtN69er+UrEkKJVtOSdiryFaOyzjhYFvvIvY0stq6ZZLL5uvWIenoZFnNslAn1FKi
kmjarFaY1TfHfK2hmDE6Iv4okUuJ8hvR/u9vW0D4ncwFvbGlxkxxIUJPAaS58Q0TZyYFZw9x6ySp
7e4mYKwCGahNHdA0pwXfyZwNj956k5xGibhzLwrNGnc6T2fB7iHtgkXPT0RwnGo+VWOUngnxZqxf
wm0Fftj4tQqtc4SEOiUOsaQoSjwyDi5+y0sbTILujlXDY3ooQusgbWx5zwRxYlrpTm6UIVYjNb6t
q/nvgDsENaeYI0XShjTM/ueC5eW9GGtySuP5xGXcmRMvO9eaKMc+OfLmhlpRofaEKXdMJ9BGNoix
O+5iY3Bimocc//2/8ZL+CdzzW0ODsErihK/JXngIX3X6sq+NUHLjPEPKP4Pm9M/YWoz2OLRBKWJL
sp/BRiOp3SjYc9k9OtUEi3qVY/Ygpz762APdiRF79e3OgqK1Rt2gxjdM1OaL232EA3ytvYSyzqKv
RnDTTk+8uGWMCZX7igEt2H4GfW+McIAM9nQSw3JDaqj8U/pGVNKJf2UuTm37NTAC2+mM/bvtNBaM
I1alaezOwT3hIVRJrE6rYM1pxQF4xL5bs9+VL7sKwLOGjQy6o75CT4q0Sb+f4V6XmlXWFcbT7Hnr
yaH3LevwRuLUJ77NlTAS3TbjuQRGrfQT37H/sDtOGYyR24wyeKl+zA+fb9iKPneZtF9zOi0A3u3t
hP6qs8H1qyhOpLs1R7o372LEFEjNUAN+fET5JIfkYaU7QBJonjU6A5dGyCoF35VFC0CxJYyEv7+n
daoJFytsWINA3c+BVpp91RFfZi9eTiN6J7gAZY7o3zHbkD3S4q5aYxJRCcMr4oDD1mR9Vl+cOfoG
CY+MDZK7EXKQ0JydTdawi9LtKfo34e8KIti5YGsktTYlVyZDv/WbDb+Zu6uo5+lh4RWtoKwJtxgs
QGmj+msItuWklnHFKG8+jWcr+cxRngA2I1Y8Vf8fR5STSdAePVXwhWMScAVQAVY0DzU/Khyruhm1
RGZNG0N680sw24JyM3Nko8iqjN3Q9Dwu3O6+PaoHRUz6IBHdIIyPTwdpLVwuuy+hvqfAoXOLVyFl
wfF33FgkvECKoFw2QkMqopwvkxCXm+vig58PnaD4nPp4DNTsK8PmmIqqq8VKp8/6F8AoZ0L2aAP9
b1K4xc4Jc150dlcO4FcsyZ+13WeG5lxZDGD11E61cokhbKkyh7T6YzpEvQpzS+zNGc6DHCrSBsqn
UTSSww5Hmg/BvFeYykh+ypxoKPDrRb2FDs80rs/mAMzPJBBytBLh76etM6908IzYqPcqZuOMtdFp
Hojj316OIgdIqzgg7yYlQ678AFyjECYuhQEupHp1JoAJ5W42rfT5kC+EVVlz6WOjN7gemgUG7syS
RWuOEpiOlubloNOt4ek8e40AgHbpKr82Ioea6fezzlaqO+ONGWTGqKCffKvmxTHCYFaONG4BxdbN
nnSFU1YicQL7vhNVlNn0bUZP/vK9mu3Bs9m68x94WM2SE6mPTSTJbICrHinmOcfL6Nx9tTR2S2tB
tRGgrf2GRSFqNn3C6lrTjG7IPPXSSP6SEreCQfdmCKVUZJ+KXTC3+CxgYeMfXXkbccn3qqcSR/PL
6bn49K1tn2d57t9CG5w8Igy6MNaaDSRuP2kVk5iVE0C38cPqmRgMshh5YsSEnY2DIJkKDFYwSFgr
/e1Xl1zflvUlf5D2Id+QYpMuvW2zGAK8SfvHiSzA4iYeEOitsUwdNljGZxiX4kF87G4UnnozNpHp
pMtCVaopuIiAQHX4DTEkCOOFt+zl4v1A8u1vpNtbr/Uu41w/6XEYFUoAJ+32Z1a5ZQ1nqHJqmnUG
NbFERU4LmzqCC6Ph8Jb5FJZpCamG185ERyflNj26NIK3b8EtYJa75LIAy+y4SJuAUZqlx8Wi8NHe
eLy0KAxsiM0CpYjqXMdeUKLMLxyoTfthT2sbJSj1bd2HeHeIPqthHYMfCuF8oNdJ29wNFK2Hp65Y
lAPR3JbDdzDx8698nhZmxsy9UkWR4m9Y7OQ+G27ywxHVBvyELnYssz9J3XuMjx+SUvtVxHfxjXD+
1K2mKV+nekvvJxpko55kOktzVDojYPWrFd4VjWu57mRGY1yQjsenLEabppm/jGQiJnx8r1sTXm+d
CZl9bFsHlOJFIMiEb+DkPj8bFZSlz2kH2XxldnwIyiKivRsY4oyPVbuM29ih1aqWsYRrJ1RPZ4HW
k6AzSLLSBg1XkfnY3n6pXg4n3vLZax5ow5W8jsfqPMBeHkpm4UY92WmzDoTDU+khq7Ua9FnGi3WY
HVYwjSCrxOyGSHcdIEhznREaia+mFEtUay+j7Egm3WvmuAkyrcVsnR/6znVD4Bz+6Tev3ZKWFVr5
pMh3GrCsquDWYO7jvA5nM4Gj2Sy6/0GdMfvwzFy3J764GOhQUd+NCkK4ILFl7dGNV3hDl9D4QTu6
mbbYdUmcHSOumbVpwXKzbBXviq/sEbEE2QULO4qXBmZYVvfLn/YjRK5XBU2tzzE8vxY/Jvl7rzTX
RjCfwkE+olbcjLrjsJasiPDYhSphOUtWdJ5pcX6QnFmnTUuN63ddvUTV/xvRt/rd8XDIjNjri/gn
7rrqea03iNlaz2XwRaHYEKyob/QMnCQj5nvbG2bivlCcLzxjJ8HaxPPPoGOpZ9797+XjOJPUlwvB
xeYlTjM3TXJ8monxWQyCAiGFNJqO9Mo2GxlXnEWMM0svH5YbMuvgdOxI+PcghJu7n16ycMVacFmI
vbOR4/LYaNAU4uFHTpzob6nnI27c1WmAHwLukgWHG46n1MRXtaAPEowyuCxG1wMYaUoi0Qo+ITDF
djIpVgbbs3kmCvstEhMR0hHgfHGh7DpUtQdt54ODycmIqO6/oTAjJuJkNlNKRVYMjCpNLobqO9Wl
YHS8Gk+f0pGm7e6h0hD6hvt6qgYNYim4bVX4igRBjgz7QKt3g8rrZUJDIl+hfa3qdyc7CTdzx3kR
xe0TsBNgQt0X81LHW5GAm2aDR4whEqCQLzwJMSoMxTwr7OYxJaggdBEgdo4AM9G5fJyLovj3P/k4
02bkI4CTDauG4/dZIJk1pIsCN36W2WCRgThzZvzljwLuB4xaDeUzAy5qzLemnjC479sERrrG/Cjl
pGJZ7eQ70D9jGmwRWlR4cprXUm5XFTO/o6NmkIml/NndQD619zKJ23FSufuR7rNA1zNpUMeHvaaG
BySixdnVeg9Cadsf9JSI1NEWRiMu1b9PekiLKOzzzZmGd2LUSf7RCiMeJmYLLqcmkZGDhZCrHySq
NYFaMWmEsEVqzs9G4th84ySwDkETKmjOTDl+DSeYEa5MPpA4UaiW9s7kEdE7hPR1qzEaeYj4fg0I
oenhDZujRsQMIEuDHZJ7ow1RdNDMah4ZiLwv3Nq/CiUUpytT/qUT/t+zmlScXw1yly62J0uDtv7j
vLOFqc4uQX56HutCmYTYcsVBa8Ow84YK4lHFX/r2wursWz9sdtzBrjsxgJ/Z/OlKsoMHZJhzgcbJ
2SRdqmVpYaGB0zsltgK0pUMDshu5rsNLVzpWmysj0XGnGaYmYyD3pRqmvu67SSGsEm3HZiSR+MqQ
/cqICx6iRa53e6JqK+sAbL/UD18C3nMAqP9wf/LuaFRbSdXQnZWmMqxLf6nODZqXWRlLNAzdBFNj
Edej4XUff+yz6UEagfiqYb7FASAOQWX3CUG8bze4x2RVtiQq9HUt4x38e1O7u8/oM/avlYilgWYr
EL/vNRcU4qVlby05cLr+sA6tfVi/W7OysmuSRfyneHvFBbT1JkifdlU6boqNt+DJy7p5y4s8p8uf
se1n7nsf4jKjEMMSkKvEbPmWI3WTAkj9XQJ9IEkCwBKmjTWVEKQU//zuLZvYPs++/tSchjqanSff
PA0LMKO7DvgElSQl0q/nQK+WZQ0580sQtu+WVrLLHX8RwRUpEqr/oL/EhpiL05DqZU7ouUmNngrg
w4nY4wYy9uuavq+Ef2JABnhAfXmu9Hkq8+f09uGd20DatlDEKSV2vUXEt01RDcM3zUMN3U6lnExJ
jlPBgFJ7+KHPq/1U3lhzQ3Il82w5CNzgosiHxLcTKecuzBlbCmWqyQ6lHjDbUsqoC9qJLKl8yxHt
4tA5wdWZuYfyPIQ5cuxKh3VB3IwZ5u2G34j2A5f8hArwX7SgGjlyH/ZyxYQfj2L/fjicspw71a3P
vORCzyCsNnSMHfpwJyh5FiQa1b5FJvuIEgNBP9BKlbgTdfmXf7w2Q+dlWdawLr50SAOcWNLu92qn
4IIptRh0crCiq+d31pxt8OlxRolfXqJdxbgB5ZGhmnwNu646lCxof8HQjDlm47XKVV2LfHzl5qNz
WP9MJmGfIZVq20hhD95+OvlYmaH1Uz8Fy2EpzSa+u81u8ldOcOYMinSDCr/7P5g/NamAqc2dhUPC
qV16clMWWX//J6vkSxzsR3gFMJYkk1l1a/vH94toTqOzqUr/UCFCUGzQwW3Q4x63bc6D8xH92Hjl
X8JMI0E036fBE4M456YnEmiw7aLQ0s2ILxXq5rdb6jpL2L+6ImNbt69mabku058A7T1+mYbScp9t
9GUwMhW9ltmUDSuNgB1Lv1k7NpMBrd5h9s2PY9WKnHH8pcieGR2UQFPoBrsX74f2IWksrUu3mDa6
qwxnRdpl0Fk8preoUwFyf0IecnM0xcsMrzkWwRdXirIohPjHaUF6z9OVAD6tZcGHXXoIWI8qwG9N
pL1pMC9RwCz1PhulzxzFIE2xjxltaqkZ+di/0nw8Gph01bPZ/JEYjUbqtfNMomlyd+ujCEfNvZZl
7+zDJ0XxIdFwpuzCxg1Fg4iVkX35RQaPdZfZmntb6m5wF2NYgZvLJlklieJwrprU4ITLsJSUxcVH
eHecTWfSH4UMhwKkoP/Km09ZEghAke0Utn1piTNQe/NCNGiZhbzFz/oCna3dmaAHeuhu9SSXbNwo
0rb4N0nrtdq6HXhwvTIQ7UrSFv6kvIpwsUZnF9ahcjEJglL6+/OqBKO89mlMBn6ftBZziss4wDiu
czRYU8Vgifwvzlmee1SvUbUHL4VnTnVjWBaeHe9RlpFvkP1dwNOeZWX/melLg2WLuINiHsnMrCfa
2KBrKY5EBMQvuezFHRoYDRFBqS8Fy7+UG82CSud2hV1/p3qiSGPOfU4j2N6CeE1LWWHQIfv1avCh
1YUmncYNf1JAebk/lcMCEJ9Udj5P4H1vBIlaDtiLyzHK8qH39GfRxiLWCCJuDxKbVzu2WGOaIPUi
Q8AH0Rb7F5wZaDehfoSlHq2jJURvDcLztIks/VLBB1yngHXs0fWU+CIia5fJ4sL3x/vugR9s6Efk
QWXmgy8KeieqkfBDE7IYR/23E81AusrGoNO46cwp2UMPU04sGBs3d/+BWMaLvg3vllAIp4Ap4wbG
MlPp4hmrB/JRGTzIeOG1/pMypuCp6X/cYs3bCd8+A/X7BDa0tcwC6hzJk3D5cPP0Mc9kZQqWHkMJ
RsiIOZiDNhcbW9HC3dmKIeTmf5E0KhBOwP0X9/IMmLbBI5bZFZhd7OW1fqBx3zPVeOuik4E4gGeJ
G0H5PX8dD7RhIDB4TEUlZwgFm3cXlmfQ/TPv0HKAGiR/hLh0uPND/H113APdTDNCruZa7cWYlH7o
xNYrHGtBjkb2i+0kWmAmqBfibKxKIN0frIKtcyff6AGdobvoBLXiaX/1nZrOAPCVtn6Cbv81O3AV
QpSJXb3vDNiK07T7lpBzFbXBQkgzx1IhtOnt3k8fkkiBFvomB1U4nviYTd58k9Ohgbcdkn3G6XZg
eb/R/Z4M5ymHEpf1XYqSrZOcSlYvUi5w7wu6cWYBgBR94VIWTaK0ENZS6tfCiP+D8B7YfhZ3/DVy
5tcKTBEl7fmBmaVojGbRV6tNCUAeA039zYAq4tg+b1E550+ndWQdM70jJt5wCV6edPC5X13UuIvM
/jNHs5e4u2jRYeyLmkk2ppvXhFzZcL/Id5NUeGYDLXj5qlVG6v9mXX2sO+z3KTI+CY4xzU4HCZ66
BerAsaeDfKuqSV0Q6o9KzWcGnMLCti5mKGzaHOGA8BwqdK8L0BYTv4jjF+Y4QS9Zoc+IqNovexq8
2Muwua4185cVQSeVC9zvYbnlrMFif1qaeJVQSvUA8cn0SZjOtO25BQEK1V6FXKP9GMrlXTYcE7Lk
/OxBOHeZBjA9wggVPMd2b4HHL9bdV5Zz+ERLm55++cv1mFPhHSA/6U8w7CjjpPefLvkhgTaD7nKP
1poCzrBVgX8vs3lwTqrwZQ68GhUpI/AKBBLI8c8rHA2nTMU0HqcoTE7GK9VoBxIE5aYAU5Mj4xFT
1szLaqFggj3+5emPtJh3iwm5980u4C41lA6V1rMxMociRAiexvFbU4HwZ8f0iyOkFgpIk16V/Ue1
qr1wNrAjA6DTbryjYK6qwwDQ3ZlWpoQakr7/7WVoXJKtCyE+qk0l2ZCPPLjcoXqzHHQppAYqdD/N
mlpPoMaBmbVPTJMGIrI0l0zDjgk+BTYmX6PZBwCcdlxk8gHHuaB9an32HT94VeSYvL8hg9JeZ5Bd
GEb0zNUsGIqeOjn1PGJhD4DMH3/eAbb+Gi/92Jztr8TxfIIwEfLR9jU7kCv4c59Trvxjo7ghyQo2
USg9cQUbG04n4CaoNeGZe/nyvldjLkABPxOy68AsWrrEzuQsAeoKMXQGPmGVQ88qYXGZGV6N712n
qMwSxW14/FKEnLLU39+DWi0dg9mwL8Ki39upo1jwl6TFHuc1geP+A8bWR5MeBldPmE7/PfABgB6G
6uG0XF7I/4seEjO5erNFfeg3UO8tYQagLoFlvD5RhQqPGRu3wVUnvHiiAYa3rKqxQ1Uv31yXpc9D
t6JKWs0KJtNnAfWA7rW39XCpCqB5ZRq1mBxdVI8my8V/3nJWM42Vc3hCAcoUmf/EMlc6wO/t/wGH
ymfbHdF/Aod27l6sd4JWcE5aLDAnuxYP5IPCxVCmVtC2jd+WQNWNyryQ0B0JENauaZwK4ItKxUOG
nkqztpv1b25VvIufG3VZKwemBB0B7nRAbQpZitFaiOwMeWuBfQgaKd3QhGEF37cFN6WbRgwYyPl1
fEfH20NKVcUuSD7gsgx6gr7pqSwITGyJchED7L5qGVxdFbQiQibtM3bitVH2vefHAHPUKD8U1SR4
4UZMdsEOn66dnGfnmpZY4qpjoI2NwIoWCw0X6aZ0P0QFFBDgbVD/xMQsS63rD87P02RLRZCq/NOA
mLU421RftE24rHorML5VsnBdMZvZQXvpre1E2t4EeAsc0XhzJogw33rF1cm8H4gxL276bJpW/zMI
2B3+Udz8zCHZAdDJM3iz2nsOzA+6bqcCYeHgC68HLjeMh54sAFTKZyPACbSJQM/DPA8Ftml/hThj
lPBoORa5OQJtGwt1r/TAhQlKNj68zQRn2FCTkiuUjojoG0Uwi7TshSUKECEb92hrrsziCqF94FMY
HE+f2W6K1UK5ANVElm1lKSGEyvRZMtj0o/gS0xhZEIiEBoolwEnyYu7bhfzrGBYmkd0untQe/mkt
COjQBaaTSurd6JDvj+ki7q6IONaHKWkg0FEtnMBzegQdjBFguNc1xQM30cdjGqtLuRhHQ8F7xBUp
D302f48Io69mysRjRkSCvMJbr25BtUySkyc5Ho/KLQUaJJuU/sDlV5rZcbrjAlYm7NtTME8vrHoM
MR5Ogcm41flzfNI/h0dS4zkqteQdu/BB20eMd1fsLhs/ysTFji39/G77kEWYqB2pf67TbyMLy/EU
mq86/W70Dn3rheQH9YBioGeOd+l3IUrWYlMNzNAO1zQkR2tHxhvILT/Td24I2+udQZl0TwGaueB6
sOEaml9V3Ybut9H5GkCIfm/UiMznydDGIshCTlFObLkKJbeRk08t2/K3s92qW2C9ivPF716xn8AO
Glf8o/izFoFOLSZDyKDNf7h3Ml0r2b9w43TIyc7hNFz30SE7dOm49nErAJ5OV68qnDNjJ9DCmuMT
6n1JzEobVWzJObRTi4Ad1BLSxfABPiYbDPK4VDdAEhhAQHc6dgtfGJzcecX6+F0BaypYDY+0sCU8
Ycl1/NhTujmRPllkYGEa+BA4i4D4tMeF179meUhdkIWPdh9h437eoBPx3D77hB8TnwsQOGIW+kbw
cq8OPIO4tIKBnJZFUaAe1gD5GGJfLCFAe14arfLEa67h073Rt0r5EESGMW4VTpyv1h+1OOBV/pYy
3jxsWmmiCXvzB49EqcUK8PpJcHmsfvvJFlSwtTyu4X/1mEAET3sDgAYvR2Q657rjA0Nnfx4p8nxo
FVgY8clmjpulgm4nTFuo5+Tyr/GJBkWM+G+BuCiwMPiKdLcuyAYIRV8YMX7eAWNpSVItW8T4eQO2
8kxI38x5Fp9Ul3NT9mLHFqWSpmHBwGxE4JTUh2IsBLkeH/57Ml95sTuWHqjV5VH2HJYzoPvYpCSa
1xHWtul4pFhUSKsOm+RZ0wfmXAzUVHY8gSUiYqWrF8L46GMyiF2zH7osF1yeFSTh+rN3RjwrrUl+
VdYLv1WWZeQfjuO/MuBNODflDDp7eONFDREIxameIUbij6iKEodnHzA+PsA96PhgLu72vta6Teu1
PdCGgBjk5Gz+UYi+LzDwmG12vfFEZmPpFtgqIIzxMGrTaJi0mhxFu42AgMF5f/Z4iCkXN66TbI9U
l366EPmOzkIDcIkw8zg7lXn0EH3IZOjcCnIKUrr7VvlN6m7lQvv7JbXcFM7xZwp5KGDx6a8isNvm
m6k50DjphpGELphBsoBc8Quxlhn/hLubzpSULNZA8SGWrv1dckTZQ0wJYcOHkOVJw4xKnKE2iqRG
J7Rov8TA2NDFPKW4zQcOvJrC22e5AJrnmFRG2jXfKxWnneIVatS1JzQTDDetvDKpDbyRncXbRD/a
WtWuAIB6ZwxK8RCQJrcmWPsbkaAXp0dZqYxUFVMyqrS0YkgTnpiLDKwyKafp6YsKfmQwq3RQ31BL
VsAg34aimW1lfSd2X1NJePLIHvwyykDBaIE1XaRmS4qunVw83O42vttqKYnn1V9EHhKd1Z416Bph
d3zUkpHZprRyyikG+BQIzDtAVW204BY9NY75/SayF83nD9ZhWss6Ph7JdEVQyCVxHmsZvw7/n2gz
JL+se8kzPW32wsjVW5f3FrVp/FTDT/oDmkKYNEaxu83nmw3c3eeg1C1fMPAEDHTF8FkQeY34S4GJ
tFLJNd5yh7ElqMimVac5TX6wJXLkNpoqu8MJtUsYztTtZTC8V90DesYebczJ3LsR9j3t/6FXaBJV
mwaaMAZUEl3zA4yw+i5IGaLa+Alid25xUQN9/rfyF2hvA1X5cD4DT7PIQjjWwsAlXWi5MwwyjFpO
iwf11M2VYmOFDgPoq6N06zfmVZusbCTPQzguVLPIx1+TrmTt791igtIwB8it6J/gj4TYuD8edXD4
zVDPDTgQ3bDtIBkSJRu0Hx1fhf9yN/ox1Fc080Zoc0l5Q7aJTUnUPFECp+9iFHeGf9B918LrdIkn
0mezvLJToR1U1fY0QMxKOpgk+zegeAm7m9sTBvH6IRbn7W+ZJ2Ji5FHp89Mi2R8GFl6CkaBaQtCR
h/8Ag2q+XS1Frldf/d+zhxT5LRnOn5HLzlc4oYpzumUzDPAk/ErhVtCMXaqgtA5R8Iwun5afi/Q2
hI61UbCrc+f79uYoavAUM91FVoYXoK1fQl7jlNgAEOnO4z2upQ4xbhHreAwcSA0Lx7bcW3/GzeiP
HmfYkgUqqtHEaL1TSiLSKjt9THkS1uYg6tiYQPyQ1z5WFo8CRqFoeER17b+3WCWEkj/DH59MVepL
BGaBQHoUKW2qwvEHaxlmryWxnzGRQA6yHdLZGx2xbibZDiQdvgpfdhBeIXXPugxG/tkVeaeFc6oq
2z0gvON4heeoQh1+PBq0fVhNZGzLo6QYhLFuyLtB5yCgWcAn9YkNX6/VkLjjkXsJCc9ZybPgZ6d1
JbyUrflhy8l7W+ZB7yx4pa1B6HDf34V/bgu2qgM+aevBAYymJc3yDl4slM0a2zwVMbkWNKB/Ii+Y
1tSq/19SBcpg/b4ceniaNtexsivQY4uF8A+XE3zk3mO0T7zpcQkJXqii0bvlS1xVNa40NpeawIcN
M5PR5rzgJytGHsJziH2OeQ86GyrRI8qxkQhaF6GY4CWuNtvMUQTNGRY9fMlFiSQFJrWXsBpq6acV
ZJxzVkNNryCrGPN4fOJhCpUrM42Ee+y8wQSjMq3E0HQLKlcbP1SX5IRIZy6rUh827dC/LMnUuSCH
pX043WkQXpvj5aC0AA4PDWayHWk2G5OTC9+TO1s2IkYQx+gxOzZ3rQA34Zxyg27I7pWNRorRwfd7
SOZepAO+YqV+YTL3wDgMFUnyf00eesmSLE+sWMSpzxiRcsLY5kbnoFzIwROuul/iBKqpGW4Esmh/
AnSMDPHnU3KWcvJmrVv1BeDtUHzvGgzooLsDS0PT/Bs6FPXYyikIZeFmDwLwRYFs6Qn7wCRiSQ2H
fa+EzywXcXqOcZjJGWhPkBBQtl0v7RBSrEyqb15G1WUZ78vXWHddMKKEsElRhvGCgjT3zGcizdiX
r7zfQKFqvtvoRkFvk4xDdAwA3BvpQPM8v0PUFLtEREZvCg7rGTfl277mjXfR4ctjEwav2YoOjAae
BNFVMUbpgc+m8gmQDe08/Bf7Ki0nKUtIk66WjdyVxkNpkbXC0UT0ViMhqNZQ7mvmKRzELgsq5dhM
l+C6NJfJlzP3x2OPknVU+SXuLqyAvVX5Yd6ozH3JBRmPx7I6zw8DNr8aBnvQ6PA+4lU0RIMpood6
iCLWKmiAHCmPIBGUbQc+GHq1IqzF9rgPrz0ScvLOD8bqIdkHD2ejwkgPDPBPbkyEhiq2ZK0Iqq5a
g80BsLA9xJm6KnsDnrklZALTEjGzI2X2nY5DAuJHZzuzdZ3rm95k33BwWuhZ5PgSU3184SID2vEV
yl/XklTb3dA5oQJd0gohHWyxz3k6TnJiV1yg+ArZ8lHkepEeYXc3spmFS7ohPllWNBjY+mEMn9H5
H3iuo4pRZDYYJYEEy51+Wbivyw38Z4crGNMMFjL1gmT7WpSPx2AOqvDSznMW+rzj1y4j0qIC7yB0
Zs4sKwzJfjdiVJulH9PC5jYDqF0Tbvs9csjxDZJbIw9SGke8HyO2WG69pQczy4lYBsERkU6/Bokt
1mjixiLegVro36C+euIgfF7CmqpEL3IjcZ5oTuTqZy2jyN/n2vIVVnoLl7dnRDDkUOHxPaM/TOtE
PnarMa+FKCzvHVSUHsf/DYG/ishloYprHNNNZZhymHtljzbU4nvZqIDHGQb+QHsWII2ipGZSgJ9H
ei9p/U4Aaymlv+rfrFv4pY13aMhHeKBm27C5mWttBQoE9gMSK86CKJXdifcPAqErbWPouv/NCkSH
uCOzJaLm1gRbQYEtrCJOo13wa4k+OvRumAcRQWDC1OTYYhdB9ZAlFcnqaKBKVVN9I0g56+2r89qe
kMf7MiISkjq5Gpi9MU+EEsC1+NiHySfIBVdOGcSMSNb/GV6dIxpHymVyxNQQkRyQ2yhC2PcBajob
LyMjtkkuCmQyCb5thUnynixoTCLRAaI819CfZb/pdtLI8BK+qlsfSOEdRDSGPNSoN3FNT2WKmjdR
By5u/3ehYEQFJuehxuqS/xy3eFZec740ch6dKll6P7jzHf4d9Vq1g2AFtqSlgT1NCgxRwj7CsLv7
L06HmS6sdtUVSFeRDVirEnybrMkOR9Vsc39OX9doWKhc8jMrYRSQDihQoU85KhuliwA9apDUK+es
QNqqfJ/nPP7jZi+j9FhExmUDZSFGCQ3jUBGrS16+d5Y67WF3UwUqMIWQkmiJqW9eOUe2YqvatcM5
OgWcntAFE4n8zHQdtUyLxT77HHk2aymYWsmkP9is4VXdv/AloiojuOU4b/cZlvVBz2ni4QDgNlMM
NRHDzGFsL8tFIMll+zk1jMoyGaPkVh8Rxy/IxYFfustSEKJ/62VldV+D4OB13gEAqY56ufuFzBur
bTcOjl12TyjqpPZf0cQ2OlSq/1TO3ulcm68HHLKnSAySBq02QoWvyJCdWnpJgbNRuynjICntTnv6
quhaA0ho9eHFnZv4i+u0zjwLeOyxyrnnfKlZsJVkXMjLTKqsNryLWyPghjMb7EgtfI3mArH0YfCo
6DrgNydnJcXUWESHvjAEoIlRK0ddHI89rkZ0jW1BlNK1gBpl6EDppHcOBIAfrKTn/NyIcpb+Ogwz
K7jihYV3iT7ECwQDQ/xv8NE6DkH0WFYfEkJLyA5edpEI9c0kr0SCEXaxwg+9WBKLdjhF2t0ECp7U
be7DAgkvAdcDl9aKBBow2kZdwnHD4IoGqCdsaNFv5P+5Uem7AM5L4Dvw0Bpk4Wmrtoru9zfVgmlD
xjbXX3AmJKircyqsuA7y3ItOLdK0Y7ir6SJcVwNrNKHPNEwV5hU7sC4oLJpEKxtqSscQosjGQuHY
HFJ5bua+rX3tXM8xXvc7rmQtuebfqBLmsn1j4x9cgRFnNnYFsbNQw6Ewurgp4eQXIafxMl6B7fxB
bAcl1N0ICleOXwosoVNK+RFdl5icGaf8PeIMmir/o0FLGRPoSc6qhnTMpXfQ1J/mLqR/6RK/KMic
stqHPX2CaP8yibFItXSHuHSKTzSJWzIwoahg9Kml1ibGpeiZAp825TiaKDCeRI3F526odNp4lFS1
w0ggvq6DLO2HMehWIlywTCmqHgIwZtC9Uf3LJ2yWIbpK9Yq9b0FRAMqV+4lHI8jfkiCCTB6farhq
A9FTKesxEfSloUbdqOsaS0pOvvgZT7ML9HgRq/EZ/tsofzMaDmQLSWdKC1hfH45sE3A9t6no2ZGu
VQOwHLk55bHVPMkXo+3q74odex4gAtAQ3h20QmowZrn2Vswfv+LjZX/uHzbXdTNk/fl0U0uTvul5
OQewtqjRtXdiYG/ePbhfbNhC1Yo6LH6wjwts9ZFYobejc2uqZnv/pi0xs2XAeivGXFqQovUoRDKb
Z5ck0CxjX0YJ9zl/iTVf8n7hgdoltYt4UxJxBiV4OH/Incot+8JwcpQURLLlO7TnIhXK4FJkcVhX
wJ6ygackT1Ho+PrMzoVDxVeTAvZUmBaJTiF+1M33CPcdyJo3S0lGZiHHrz8lSiB02Kit9mfQjrMn
Y+hyVFyscS7a72oaG32kQpftyhMBK3Ic6uIKxO8ZbfYGhUEA1pzPAjsEHAkdXVH1UgxTH9HBpkI+
6RDjqOv3tx5KHcU1VuxuB2EAxoC7lDUE12ZS0a44Ct5EpWuSqJuQRiGoz910InDiLq0pwUQ9+m5x
gUKagTctn1ahb1pk81W5MaJAbXmQNnusGGUbSaXs/jkLwhyQBHtaKnY/EXBAQNXWjwXpeo5gsref
18LJ2cH915ji3W2dmfifnvHkh1AOfS90ftnj+IgZyUiHjnXEonMYvNPusI93+5MtY6RhlZmIi91H
GH20y9VcPDDSn/tXmA1RTwrJT+b0VMTdvOBrKe2inxg4yi9h2Q/I1yvxKHEgiibr6DNiio6F8mYd
nRhtgkCF9pXpllvCin0EOKB+4LEQOzxL8phZ+d9gOUdB/LWs9tJ6GQfI9NYEJtHfr4dzYz9wh1hG
N9I+RZYYHWwvTkg6APd4H3knQVvi3moJeoMJCxLzrAsy7cFVMn5hNp2wv6B1Xcep2F77VeCx8fMm
eVONTPWCzylPTx+/VHqFSVp8d/oxyfPz0qtFXIE0frLEV04efUnj8+05ZdVbZ9pAaBaemz75nrnW
y2k5Ez5jC8ZScmQnOqgZOLSIeyz8blcVSj7fEdVeRPA6RybdwtevabfoGd2OB14jvmMh5CCTZlrx
ML3cAjc+Zvh7i62FE2mkmtLYBlcLl286B94EuOecUCLxg3Ci4jYfWe/YJfksjWpuwMJz9k9FmWZv
7AZv/OnlAsLMT+dZeTK5lEQJXO5FmNKcJ2ha/sNfCOVBhmZ0OYJjhImrp+wkz/E/jlymc1wlLub2
BqmxbztNEql63RHjSZv+tM/I9Cf+R/crsEKD0HyxjROHU7Z6ieAutisRvWM5tUm0W0bLhlaRw1EY
v7d7lLYwVqsfaxQU6bInzOZHJlJsglI57uaWi6ibwQ5g29n6L3IL3UNz45B6PdT7mqJ3Vr1GlAql
otNXfZh8PhyvrEyp3uVp9H4TagwZK++P1NSYNbcnL2NfpoHGEsl+/w7g8oOOhugTACg4tZYFY2Oc
OYRLDQxk1ciF188qfp4/yQy3YOV/nJ8vNIDHo5AtnweWfYhsF4zttzOFE++wwtQSycltM5P6+Zz5
LtFmnSI7i6EPv3guRcpBaXdd89edAYXfIR3qbeOd4EiFK2p7y/x4oACeTVKfkvfiSXLWOdj2786y
XG77s6RR0AqLOrmlv8fngjsg1dTQzHVRQTx05oB7+66uYYO41skgVDlamHfJQBmuhmyoympt9606
u1LV7h8+torMe+FZNntW2OCBO16oc7+yEVkBScSYG7f0I56qKgJMyJZGR2Ka4Fkc3zPsMCI0nFdE
off3IF5BvFpGowt7Rjyqi56lG4XPEmkkEP/KnqgtBYyk2JvqEw8nOelDzzjTywctPtfr5qzFFmdT
+pWYBlz3A3tGbj/TMhd/uShQqK/+/ZwKqfMxFF4ciS7HcjO8CWAgwQm8PTC9umuJZCdqcl2yqU1r
zehO84SPWdChxDjQyg5g6Aq2bQryF3TJJSJpeA2s0bw7byufhHqIVzhzUFIeR+kWLq7PTh5YSGPc
SFr/J50hoTCsvRheAXmECXWiOHs9spM/BxiKQqVfL26iz+Rzlthr2cRtVlVBnO/E7MxpQvlFIDO5
Kj6WfXPyl+rNkXyt7vU+c02HI3sPREqbpLPVvPSjAJQABHdzk1zvQ6Tf2rd/bZt+0cyhxK4U5IDd
GgGgEXaH9w9CDqB11kYglJx+Me5CE2r5l9o0V5tO1fFlvEKd9/4EWZAdaW1mQ/IpUf4QYOO0LaXM
hWNUBjPavfjJo97ud9Qdl5m2tbpvQxHIVibEnyaXDAuqhj6KFrgqiR1IDPYlU81i0vsN1kO+G8ni
r82IfcbzvBk+sE4rRf5vsHmBC7LmurxsrezaDEHhTnuGtOCLcnCoSee9DsBzMXJbdbxGNZGP/Za8
iXMcBJXVyrv4cbtzeDSGp9EkEDDk3xikWqI5vvuwELRpkxRXFIZ5rL6fi6swRLYOkIfTapWyr1bm
g3Z5EleXk22m+CEUGFXKHKi1HI32vSCqYk4D6aN84pn20Lz0FTTEyPDPzgq+sgEyn6jcKxQR1acR
ocKcwM5egL1pAdI+taEQxGXOCXs5PiCz0tCPZ9vTqb5fv/+x/a/HY+l88Kufn/66NcTQRKG/eYIp
S5AO6vyzFoYug4et7b2iIteKp/jd/f0l0o6c2/kFjPv/SIxth+aAxEEwm14yxVtwzmxlUuv+6P0r
fRTjPGJufQfl0osH+AAWiXuMPqQyiiUGemx+s57eNP0obq7HlAoSaaYsxL5Xbj2RqqYGWnmDucqm
OsayXTJPQrZVdt15rGUmwu0dUYCLW9lHcCvDyLC9Lxf895M39J2zJVbB5YuAN9CTr/chKljKL/B8
nOfXq1v8rN1N9B8zaub0GIizKm5JoLlLbcDYYgLNO0wqGf5N576WtRb3KibQ3uW8ZMEhe+38t7re
iIKz/AhN7ljohEBeMzUkkPaJh+Cx+G2C/nJIuoGSHh+Lj5FQudAXtnk2+a3r9OZVaJpxXNx1gJLQ
MDzq9ZEh7FtLdF3i71B79u+RttD/R51FWS2P0Vt0GVv0DYzNt5i+Eo+eOk6RQ1s412vfFj+duJmo
JlTBWlPE+H/2cDmGZQ5amtFVey9LBBt6JV0h3Fn94e1SIH5EhKj6YRqFmzaHb2xzK0SXjnxXNErU
WtTnINNMcUyslx5RTYTfR0PoWxkWNqMFMj7iz32Ij7SJG2XImTKwRGLOmAaOalJBURT/8DJYH9sA
YUUwrCjT6pA+91cRldB4yKXYiUlB3aKUIxZxWctWPxkOaRueNjVSAD+/7nCP4+laCC+IvTnHw/u4
TmMqdrwr1fHoNzotwXSQbykzjV8eZ0GjbGXQzGZ2AY//Q0ixh6vgB5ldkLCPGXmJqA2ajPx4JpwG
lXar9bnjzMbdAVqvJ8GrCfsjeYl5XdQyaiCqu0BgvrWFwwq6EDVwyCmjVD57NeEMNkPi3C/UjfeA
89z4PLazotyfnm3VsWJCvNyaI6QKELL2fKKYwUxjTl1RUjBqFN5ZbRN/woTgDeMyRUG3cEIotRPi
5prw20KESl9NMn9hLzw83pEAeVc2+tYsZqjZhH7idrD7vcxeQbrOE/tKzyfesp8gqkBbTWSvoTME
PxY2SgQC6DHwU1vsD6i2pfNueWLK6tDxvGGDKjCmc3O0745KCkelFhV/uSgaZA6Revg3Giu2QRXq
C+K2pLLY7hKh0+OqDYT7+w+ou+wScUrivTjIW9f09F7BwNOaIrhPDToZC29eGRS1XMm45hnPEm1b
5ItiltJNIz6GR1rx2aFJs+8F2wDrjTPQIZ9Hr8tZNmi7uE+dcmO2kVFs3kk2YZNTy0aluc5aolHV
qJOQ+eXxmEs6mf4t9/34MF4OAoss1p96Dm/LOT8OIQjCnBBdyiyD7vEMGDEftcasB3ZOEKj++jpr
bovuyNOyrfJ9HS2JzUnprHWkRIeloQ2y7bn5DOEP0j6zkOpL2Bsreu+9VwzDEM5l7hUg5rlfzIie
8A+dhetzDSAL0FLsPRMsAuRtXQp9ouAnWtAOOGm8cbpJpClC0Ryzh7oztNVdfKDq7qRSUSPtZrh5
oYxSrN/y6kE06/K64VgiMDgeWc4K/Pzp+xvAsQukaolokFEHCZ8JeG7sEJIkq6YDBh6/YUbbcwwk
AVW3CCoh/8Bm0GqKJvGfwKY2GB8MDh6ecV25ke3UV4dXE2qDbF3rt+ee84ySh0e35j5bjEkgG/gv
of6SE+ZRIUVmbzluhPDbfWf3jJFG5D09oB+rlrSX0niEwu3FMSRURN+0if2A9NqRTSLiIsi/mOgQ
GUSlCcGZHbXdMzx4ITFvZHLXV1XlTMam/NqNldoTa6MZWPOnQwr+8czyBGpFNXr4hZsLuSzCnW8X
82oP6gUz+M+N2MXt0x8LxIKPfbSQt0HgzX/sgPPD1uB9Iyy4s6vt/yxq+0wRjXqEk9yJ2ouA8zNC
Ihg7XWR/+AoQoL1qJQHMEywIchLZNl9RA46ZpaG9RavfVwj0xVuXDlDuylk4ukxpusFFzo2XyU+t
1rnDE9P61xXZ2+SGYqCSxNfX+4+f6ICYaDWfLRUfRwFyB93v5EBY0r+xDsaUV0FIrf6+UMi+Tpmj
Rv/12nUQtnPdw7JYanfq3x049cBqtVZm/pQM6Qchc2vVPAcdGtBKcO3/d1GnKQaALtwZr9nK5K79
ZRri2nxkqefpnVdkRn/V8eblcqtitqbYWbiwyyRILhQ1iGnfxmWcp7XkEWYanhOUmgDgxCXyMXp9
ziDhw8rD5PL7iMNjbW6C7Dr1QbrQMWUhzcTvj+VgpCw2/bWol9Y5f3f3kFC1Zq1/KlETdjxVFHu0
BrVw2QVVcedwO5+kp513e/38NzBmW79+9RrYFKIvQ2+W7AkUWBWn43gauxi4PPacUjEKNe+7Zg4U
1ePj18lkzlGxY7UVcq2S0mSJ4SKPjk4DMnz5dRn7Nne14OSEnvcB5JEsiJF7k6iZ4My7dbaEuVTt
52yw50IOi2Zn+x3gJLLaN6aLWIoW3Okf92RsdEiSwGXlF2r3N8eHGJS1i59rYPBhnHBjIEo6hYYm
rYwl+xW8FubM24yHrgxyFOTIPzx6Pc8Kl4+alrkC6D42sV4085zeufOdS+9eteRpkQcoe6R1Imf0
hK0vYfyNPOYEFwWIkZWoQsuQih/UXTb6fENkPNliVa9UwveDRl9NB4ftqNjHZPjGq0bTCMkrxJx6
y32uCmXQ3mDkp6r+mFLzF9D3mTPgoWX3IeMJJBNPKzhrpI6BhSo872H8Jdkswt+v63L7oLwmjm+K
SyDoxz7qqZKIgrSPZsgh7wXyi1krLucUJFC2LjPPmGpsJ1+/Kaou5UYECCG/BAHSFNrvmJpILpEV
R0GuO5MZTjbyt7pIDWzUHfjuRiSKox+WZpWjvFpNi1KWgPh46KX5m8QLpLCZ9dKFrZRUEogM0Gbg
V2KITXRzsHqDk/DlTNhU5zxrCz82407TtNwcb+rphHGJ1u0TQwfxqIXCKHkJcWlS3tMdscQ4A84L
JCza12QFE5WliLsDwjMqmyJbqhXYdd+5mBQvNreU9h/fJbAr6KeglOTYaDMYebYCO+ALQnvCZmz3
nge3qoIwhpa2Cm3vgzTwQ53W50F3D9ex4UPNAbxLEhI3dZytXTYoGHOAlxG17tVQZS8ag4UQGW1B
MCy/jTtV2SgVt1zboI3tx69eAnI8dr4c5KjJ0HtlsdiIw7FOrUVuPz3ANTWcmathN6TL2WSmQBR4
XNI9/6WFYV+wZH8Cieb48JyRQx1LU8okX9rS6+72VZsz5xKZ6cisIbaACsTFg00K0e0GAmiwaGdy
+wR5/OJbnxLufJltRku7W9uNN/oUGcz+KQZBZcu+vxjVhi5oRsPvq86QFOkjcGwI+5ASztsxPtSB
42Y30Wx1dcoI0VxS0xR663pIemx5z0lxTs6qIi0mfW0sJ5zx2m391/qWC2EGWrjpzWENGHSLx1pC
ez+kKTVB/o2304uty3mUpIH7n3zo8AufD9DIiNN7a9QbXL7Snf1Lrcp2SObRkTJU/qOlpOLSgtsl
nFpOQvL4Q0HHCyS264s1zIN7jVjwFkRJccFLO5rBLZKALIOQm730u3YVkEH8pfClLmfMBdPrQRM+
ve6kOOeiriGLimsMVPFIvnQg98Q4Q/3i/DcAqcIDi/0I5SPoNbK+Nf75i39LfDN8miyZJ8JKX1I6
tEOSZvTfULb+ldfhh6w7D6LkkgpO20rykOb6i9p2U0zRvkS74vwrgE80CLkcFbrABcW6mM3rS4zB
wdNlipTbe7VlxfDYptnSy2WrU91xs+Sfr9Z3q17PosK8XVvqlGAup5ewYXAVicmUj+/9Z1zu0Dz4
BKKrbJp0yZIYDNn64orL/xEbhPr4btOS8YzIfNrPZ/OQE4/T3AJGoH550ATgZhOI5CH3jCGgm8zY
Z+Tu2LfSu2ewkzSca69OaZLdoY+avqBUFO5eLjdsIFMvo6AP74XUFR9cYAq0u4F0EvCondvNmMug
2x8AiH5L3VWVTb7VW1U5dm8EwYBnFMkTokMIrAgPO9E71x3IYPbYjw8XAeYOs6rZxw3wsDA8exs3
ZZdeiReUhq5w1xJDF7+V6EWEGHLkozJDbL8GEY9dIUpW5loo7CnyYHIRiPBxZJRR0UOOJCBmo7JS
mHfayUyWigQC4J4bb/Odf4VXPJpG2fbkopaMvydFOxO3qxInWV8oTcX4O/GK11U1OYFsAsNMGGGK
osDeWrX1otGJpXyazamIIuejAAQtDPA0StJBRjDqZtvqVFxEwojFdQ81PsbHhzUX9+Jom5mJslo5
9CUmaYUn4ZrMGc5OdCERHnh8YN7fOyPb30dHsz6Bj75ntacIOnkcZ7bot8WC0pFIqu4TEW4/59U5
/izD5tplnWsMNYOlsTd9MBbkfbhrrF/rbAZAykl/ea8Owb4WuHb7OwGkYoePA2TpOCPJOqX/dPrG
oZh496zaR+91Z/cAx9MPXUXL7GK1iA8mStCkLwm8m0q1rovWT7A35ocgK59ToMk1lyKItXc1lNvr
KMFrrWOSXNYkdRGCIq4Y0Y4OiQJ1bsaiLQmNxBDTJdEvyoxr8gx6k0znKFMkL2unnf/959hswn2U
Vv74fSeD2XpyRvxpMOidCTF4Bqzte/NxVt7/wVeRH8sJYk27okzz/wqqkLG9xfWLtfjBRAHAZI5/
gI8mWbMqzAcOQTNDmmjHlGfZkthT3MFG4NoxP6HhfiaFyNvlEx4cwbk1b//8XCSC+CVnzlL+ganL
upFlCBwx+VwwLGLMBrbgY+M129fwOUdkHGe9Ye2Qfc4XgLywXpQheVPq5CagCG5JXeSSVv4hte0D
S1ThdMrMIR5Yk3E03AjZNGZOJFnUPNbVpWSwody0zmAmOP3hiXuF0RFxQCJFdW4cmdWsGMXtecus
jd2/RV0l/tWgHV3tagW9FUY4FU/5JLGSl/UfnKZ9IknUJr2lIYwFRd0gAVX9XFNTo6FgXH0ff4WL
h19Ami+BwS/EJYHNo1vRCE5aUoRGFC/Ec+cyhwLs+TItNe3QIaDyUeIhWIDPOFYZBUBYGsRMYPR5
V8CigomCY5lBX6Ut6hjv1Fdm3nC4e/bRQa4JrZk9Kb7OkdrTdjAO6J00xTZxDUISPQJgMz8waeZK
ftPTgXmbHt+928KVB19bV6eHKsLAu7wSZ9t3e2qy9efcfND+xkBZqCgjWgaRgdDocbiYXv93hMMu
gZTMq9JgXveE+eRzmsJ5xgXMC3vVcEFF8UBL7c76CTEp634NC0lgddAgykzHuns5vYOYSViSx5e3
m9IJGzJEl95XvpAF9bFbuZG5+c/LvzzTCVNG8Q2Aj37vpde3mqUNS6dlfWcLyPsQ5oCa6lUB/DQH
+ScBBbzFyy2uR+TrFRtXmrjTDjLPF7SmWaHu8PEIWBnz6mEk9ZOg4MSJH9D2nD7rYQwbnEWHfH1B
U7R5eCMqvtC1VPw/fRzoQn5L9m3H74w7INP15vK/gvwpTKAFGCEb4YDGz3A1IqA2mj8YY+mABuUo
Wg6g7fPIqKiCgjTDHS2EB0X+Y4ynwbe4SgVMBEtjE4kdfezuHX5J/JrbVL/3KhAEqBc4sLocTsJy
TXWzhwW5DelmuCT3p4RsXIL3ZpORdto5jYc3dieQMPAQkOd9Q3q5A5rztORpVyKFd/LiD/5PWK9O
PpW33npp35CFoyNR+5yjS3u2tY88IO5Ygg0Y1vzeFoXdbOwBjtW3Ue+EkCbrfENcAb2V1Zld2udB
bJIbKQfAKtVb296KHByl5UIJ55Nqyavu1iMstOu5054QsTRlBtHAKzKHLPDsl871/Zhfk82iHt0S
0eOqpybMm44G62lvrxFtApzapUqH00i936EpBs1wjmm4Oavbm3QuMLT7V7cjT5fWcT0hNY7pIpQE
vrPoQvgAhcZycHNETRSUuQxdNocIuOpQ4SPPa3RjZQFahDS2vVWl0fLUfLkMwlvnpSN55JzQo2HS
dySJ6eC2J1kQqTRLWBTSe/H1k/CXT6ErFo5oCgNFjCf55GLNricgikqDhB0qXUy/L741MUNn7yu5
5ISO3RytsmjUqMQFNS9lJvm29dPWGlwc6H6mtZG3VG2BFJn2hFUb97rU3lsONIofozzWsMPVy5qP
sHneh9PfvrP1wdDo0l1zmUsMu2ZwsrqSe9qHDM32Oznweyvhgwt2ISHh8DZLbx9CnDU/5LymKXWW
NgNIwt3YOdftzFqzyADhaWZMSMuhkC9WTK2WAmuhUYkJsQk2r+Ufaw9BUpy534S5aottGLUHfdQn
hVyuomXDT6FfF7+XJekVAgJ9TaB+ee4tG8/k2yAEPmuqBlUOTOuRuDH7xQLqMCG1zs+CqToOQDNz
5dfowxD5mE//XvNf5ObGSxKW0DTcYk3CwdMVG/G1PYcFUI1LaDC5gA0VW36nIYpeK/McVibCNqGm
NetSL8ogqGZv1S40CWeQjIcfGD18B74hzt0BxuhR/AHLCrBeTs8Vjmz66sx44zBEDZPJEt4OWRvk
BqNQ8ppAyWfF7pQ7H05OZL9K/AxVadHwFpjKhRskvoVsLiATcTDF+ktPTbijjluOyQ++l3jBfOa8
LIPaSsMrpdC06AGXTaFODHOXenauxExq613MP/7atNgsg1ToBgeCCFUg8MtJblCxa41GHWsV6Wqt
vpyIxMFwz8JL1zZoIo/qgT5QEdf+atY6zhvAX9YsUYW8MOdWM3J/9M48NNWIgfil1hz/hNyOsQdi
twGG93gLMYjuVLi+Eu4wdYMQFJ5FcoGTMu8k+cRkEOQeheleLlzKMwraOzpduGjMB63qyBEcQuvM
CI/jNookuPgSY4w8jNQFcFFJJ1SzgT9cbapxn4UBMpK76zeon5753OFHiXNaPrIccLMA/iADmmgJ
oakb5S/2z6jI17WsCYe1SbnlktEFfuD0rQPhDfGzH8px4abgpd9k9SYusJf4M7kg1DS8NYpzv+6E
0FXF/CPAbpP9OyrYZuIflPa3n+0Ts2UxEK103Ych17yHGt6DH0bJnxWUc8xxsstg4oQBYvTXIDlj
BYbkv7wiwSJxufCkHsKsAcjUbJxgPy8hnhD22PLGAomd889lNdaHY+g3ib0KOsg3sXCOwjvmC3K8
KBXDdik7gmv5BzXBP3qcLCjmEEjrwwBMTvK6H1MmcxHGMObv/aisfZxvxoq3HvNnj0EVCp9skYPP
pW/unTrHB56wZZmHCj2zuCeDpelcMADrtq0ELPYhKma8CZwftOh9hBcMf87HHJ/NhevPXlV/QlTy
ZDd889Mln1nuW5XfvUt8hGeeQAyQlIQsrt9t5aHffOLmdhQmGTN2ucxEph/wb2XP7qGrNp8IWe5/
+JEEShJCVOTAaOuDu9PDjvaXyB2hu3bfUCAs2YnsGWOfdyZP5mBOolqiNuuoipci+DFyy7G4RlgO
glou0KkUZllhf0XRv/TS73V4wINZj2yPeEzrtMlnmPeg7aJpW5MdwRZ2mRNMCohJcKWrV2omr0+B
vuBtyA/HsnnqmGSeiP8A2k4JsHRblfJJHbYCJp8gL+PI4mn7lU06qKy1kSvFwF7uqz2QfNU1WjAj
qFW0S84xA2Ix+Nv+1N94lK/KgGDwdnZtiRL2MeYz2ggIXYRsn9swYNTLjesYDreebo9jW/S35SFm
eMk/+SkE2xrlF2jN6udgacFBxtszI23nWRehv9+ZrFX8HxdCr2zfLVd0POxkvLETs1gb4h8/7+HS
+5KWLD3uOh9pWzy9Y204p8bym6tsrRhL+aeXBOq4kxgopg89syvYHkSuiPAnr+pL/ek9sh8Q9I91
2qjOZdMW3V57UEoUxn4Nhb9E5thNjjXNjMrXVP/wLToHGjGXzWC6h0cRJivUr3Az5ADrlh+zSpTs
4r2rWPlthE8ZxotOmgYs8CmYmWczcxp1yNHqbkqFfKpjSo2R4ZySfSuXO/zMH/43Uvy5kIbjOiAA
TDpiE7su+q9o2VpMH809+VDdNKQOSI3ILL0C+XLz7cKmbOyr0LrTH1nAsngfNjFhXhIIr5CSSD4c
2wjjb1tit/eukhdlW3Z+GF71C4hSmr72GTPGLWR8SOG1aSJv1RsJ4SMBuPmrBA8g/RIHtulgO2eB
nDHywMTMcgQMDRrfGiRxXY36EGG9bxPn65lVyTE/2IdUijK5J8MZNVWbfx5Dt0kIeVuQz2R37DLe
qwgotiw45SeVYAbiTlN1T8VU53kx6KGSo/PKgK1glNjPQzwlu1y58HxUSkzdySdGXxZqQJyr8x1+
IPLRK5HvyEq4icyS7+yCR4eIqeuZ9Ntx2zhk4XrQFMhWXChGmqwUioY7CL6jtEBuY0rBod11/MJJ
sfmUz5/Pn0aJHeDSp3VEpT3hu5gAukZwMOcxtKkj0ACTq+tEPdQfh9vvtRtU81bFl8RiX0FJMASZ
aoaRORpbRx5Bz4h19FEByhhLb+KbSCfXfIR8BWCgB9Eig7WvCoe1Y/bvVrahthW6cm2jdm+UvOlX
+3403pGKJh0NqVPJF2TwGOxzIKmF5GMCmXupHxenj8bigYjBv47lWVj8o1wdEHkB1DDYjBBRx6xp
/uqJ15kapsOmEMpFK2o2U0QKKXUHYYGLJ4AOoOntf8i2WHdPwsRF5Y+tjdVxiQfQ5Abs0BHy+ijh
HBW4rxV6/yHX2J6jPRjVUC01cLaOtl5PdxvpPjQKrhEAm80u8wfAC/r2GbdUNU1eDbbvQ/x+/GgD
B6MhobtNPsY3nfDbcBQt+nUucXLMTDyyjbb3H5dFNTGVN0TCOFzeqGjSvDPkH/kqGj/IhIFLGJ1b
JVuBy8VXIpZfaenoPDctXUZM7ubAo5lHbceOCbc/0qOJs3NCGxvtqvWTUAHjDo8GzSD7h1hCzNB8
7M7JkB0BtJ4ah19tePi8F3JTMMDYvCwrVKRXF5mm5tvtzeLxJ4zwXXwjZRTigr9IFqTcqyR28JwW
oYF0LDVkLZVsSuKhlJk4lSP6XXjCVXvAH9c41gf7WMRtdSgUzyNReW2CJ+P8G5hQAz24mxotS5sW
rtfHUT1ItmVPhR4MLrAVZsdthPt2+IbIpWrdPlXl5924Rui67Fnu8wwf4sb0E7K8f+Y/Vq2Ecpf0
DoOPp0AOB90gl3OWsOLxGgwNZqDZQjYNe8wteXlozHP1klr7Z+xcPvX4ifJUHgjfcdsYt9ehNdmI
51DUHxdlmZLvfTxfjy/JFLtNZ81H3kMFRQJoAa38jyMzROLTWoTAgSY3q5iGyyvoMYvjj/ogUbGB
D20NEIrl3GmzWZybJaYMLLWlrx53CFWMA0vJdGrzh04PXHnUJAWdMl8pdtZi05WIPZ6WpbNkoZ8w
BVtlD5uLDGvvJ9958qYxV0Nn6hZYXgqYjIkpb45vu87iFwuSMfRCraRYYiVk4v4UCQzPFTgdPW15
Ly8JqS1gRHd0Rnii6z8u8mEQXtGkHHI7LS1wAv6YtiPIuJ8kysojQasV0/AoIKjbYnEF1uj46MCg
bbwtOUJ7jGqRv5AIITUBN/ccBj+GJySVAyBaLGqLGx0zYQtPiGE+EFmJTwk45IXXNcuhir0CNd6p
26CB+7aqOb1Oec0XndmoTyKt1h6ori6lYiTyOACURk6+8NRY0RK+n73U7KhfOaody8TjWLBKbT1J
bhJgPFYtcdoOPIiZjc9B3qWxujlzSCin5jH6RKy7pJaMyKRsuhUtmuS+79InaoJGE7ZgVc/1GZBk
Wnb+qTQJWuU1ORpWjG/DZpdanm0NLb18FNplxFUtPaE1clxrXxzB7pe6ngwkf9JgZdBPH0U1OGbH
d9+Gd9jnOFXnKc8sq0p8ObrHqVSX08w/voAAS/u7YngTOpZYMiSWzdWpIzbGihlNidpIhFQnHm30
HiHhjal7fx2f+OVpJp0Rd5zC01sB05l+xUjsPKKOLTGxY9xawb5WMfLgRkzTR27ttznjYOdInX3b
O/KhyjtWCDj/eDV3WBWG9npdD3xngeaHVU9vHsgeQMqRDdOqIsnITPx6bsqn/I3hkM7Xw97I+JFU
nYBTbuuhNR6P2UoxTd1w73tPpoTd4buEnobP/0E/SfmEDZ54jcIhv94XulJeYQXBlG4f0NjNQB3w
Njflw6X+oUJLZjfwS50aM+rAvxiMWp+S2b75E7zidbXCSE6+M2AJKVJRKErYAZN4Zr0KRUSAIVOO
kFD679eyPG6Zfwr0/u9YhujBxy2nu1kV6OJ/P4ciNhRmGZCsEf96LryzB868WmHVx/NQ0cfRi448
dJ7fzzlCgHOhgzpDyBGr26Lz7UuzkNG78Mr98U+2Bs1NAlpFw7DLRBkeXy8iNe07tkTq8yPivPrg
KkaKVhsq3zGIWPs9345QMbSrpyZ66QccMRPGKahsPI9fZk8jCbo0MHSz0ng9Gu6p16RuIDGoGQz7
8DBj4dRC7QVWUL5074JHQOfxTBiu+bQaPlFhKlbeomadty/URxOLp5OPpdOzPooLNUV39AXsrvEx
qLg44zuHhuff3ibJd8dVsHYCKcN5qNZV60b8Lc6abBuc/+Mu0O/N8bpkuSbyEM3g9F34wUP6vd4n
TBtKKRc9A3tCGSHMEv0nVyVukHZZhyquxYmrGQk+C6pFHi786ri0mmKL0CRHvMdywiej+Y8lqyIm
IuWx6w86+41jtx2Zr2qEKDTHGn15s6ULHcASgTGypUAoEW3XsvKlHR22vnxJSnLjbHiHUScyZNOt
jmF/UZ0gZged0RQ8agiuA9mwIlHM/qEyplUGONilDt+yidZJ3xJOP0x1aDjxvc06iNMjdJEcOJo8
olN5hPeVhQeHS6xZlkzlOMNT3WTzGdkhh98l1V8pmmxfhwhtFsPMwXYM+RI6Y4mD6h4zoNY2rhON
6H/ialkReR716DCtCbNl4sfVl64lxaleplGANS1AW9NgqncykTPhqGIIeKjuj+dyJlQQ7LrOtl0R
sVEOWenhmtZVVEWzjqKnGK8Wds8DAU0kZAWaoP7FuQWpStbTWxDm59De4iQW7/r82vVBkRy2eLT+
c1sQYqusPgjKSVPXMxF64p1ATjrJEBMBqFIb2RjvUaCxhLSQJQrYLn1wRHNVw/ZLae1F6qQZ9Ws0
AfQrBSyrnptdABm1xJKP/mc8KslRwWkufYUoN7P2k3OqiM3uQfFL1VyxMw4NmEw+bAU1J/QxRSZw
8EgFkkQ9Tzb4CMwwPJ2Zb1Pt3We8BNyM/Cgn/v+7teyFCVNBiqzVCkVb4mS4//C4fh+KXX0FWeVx
zsI7xZQ+cPesYCsnJ/a2cNg5GOZEdfa5qP91MiOthOSvMrMYKN9OtBRj8SAqwNJaINP9AfdyUeOf
KeyiWFj16/ON5LdCm8q4A7rMDbyo41StQpCXiU0vNtIGg33Njdvjh8lgsUEO1NUqpwEq4wVxYp83
R/2FrVYUEmIwuRir9tXh1nzCyJHMGhM/8GdqF5YcfPHJfoFH7M9Wei6uk6NLk/8mOtVPXw3SHcZY
8Wur6zwkjb/LQYK+c1X9VKgeoz3TbAgzUHFxAAsZ+XM9U1LvMpydo/ZPljo9iMrEx8UsSydg+MmB
iMCL6TBhVw0CNuOaHTxQyPQ1WHvZIGroCKsniKnYu8KONxXohoKcVkR1uowtfjDdb4LCnx+fa0BD
CVK0IuyDVNExZ1Y9JjVP4n1eXbS8eYdBD6xOQXiv52QRh6Lq8oHpYOUoIgeK9c0bV4gHE3irQRQ1
eqH3BXp6f7CJNshQA3OZStFNDF8Ydh3eIynVZrgg1bZTpJ5xPspOU+tPt6LIRShGWSpRIVSrk93X
E4SM2BZWaa5v5hyDa9HfZShM+LB2nsdh/LFPR/Z919OqZXEmhnsAFQNE79HBDwLH6Z3pVnd8BvxO
K6muuhVVC0Ezjup4RuSNz9/gm+Vfsdb4L1mRvvplbXq6OGtz1EvlNSg++6UKmceE74M1UvOSeSJ0
mf1Av7nwrgDuopaiHrphO0+GP8u0ZirXQwxTUKPjBkjo41Gx35tYyPaZUWvUvRoVe4uUv6SAFAiX
D44Z559CW5138mdoxgYIFplvXdIrirdfaDNIx07ClYMZLUZ/ur5cPAAU4WWbNZ4Zt0HUKUIAielB
m9dafbyHdTzDZh994Z9+5lKUVDSl6gKPnp9svkN3nHa13o2L/MBEVRcLv3Pdk8W67Dls48cIadEt
Qb8sLYr5UyvtE3LZFb+ATizOTrU4YoI3hYDIHnpkZ4Ecrsu0+VPK6R0aA2X/IZpBOllsqiw2UWaa
+l68wLrlkwdaSb64lNkx3AXVLeMHg/t+dVXXwadVOqP8SLiUMWV4suKhbLbVVi5Ns8vquUbQVXAX
uWoMnfhOvbc2SETWvk/7OOX346Yiwdba/BVlhtJZ3sODkOQLXx84jrb9rnkkoaMpt12TSD/VD1fm
Oe/+vd7+0zk0uWSRTINWMDjTLAJkGeVBldJfJbDAWxTjM8HyuQEZ4DB4WZGF+u6vQXqhJhi8No13
c5WKdHGNDcxC1lEyQa3drdlPvG1Ssh5bx5HHYN+pc14rL8OWqSnNaVsoZ/KC0dfVdAbIJs0UpmeS
yO2oJ58pHcV7Y79PknOarc55K7WJUjjBPe+CraLW4q2RPGG2ZEb5fQPmrk75kgdqsO31KRnlgw79
nQ2jNx6wWkTctdK8OEpeUv1IoxYIn60YEYGBBAowkaVXsc5sCzE3iVW16vhfE9SvjymOkeAzTuDZ
qPXAltKiK7oJ++jap9VF9joEfm0F6WKirJ+FLVbStnl5CARixgzZ06BBPL2euVOvyQD86Nqn4yzn
24kWyLieDIfIwugKtWgBoYKojGdXO4mWipwHfnHZHip+WDtoZ8Jl5qlRTNJpNOSVCndA5C/CTyai
nQz8e7lUOKP5zMAywVXaKPQjTboyfFt2WiyERwhv9f+UUrfzoe3q21Ii4zc3L0WZCLtY1IZOBVY9
FS3F8l388Wepbs+9NxnAFcddi4rep6L6q9A1Duk4t20lTe7SqG0hS5UCjlMjnOeWVbpz4GNQs3vF
wD2bQq8BL2zlWdxDRD/ls8z0O2oVjvPxq/vqscvBiNNW9ZlhObhFaxIelL6M3YVPDyLyMQUfSL1u
RRynk2Oih/YvDxBAiUJXMig1Vbw28JWKVRCW+qMPW7TqVB0fVpCpk7IreAexBt40rxIOs7ZEegS7
/hoUOwnhfjDYjhOrTP9OYhRf08/fanUu5q1o5MFRvrCU2tovfFmCjiqLlRq2CW9L/PzJYn5Vn2wS
uLdB0Xi+XG8l0Xfv9f84FfBhlDehbqTLQ7q/jBQ/iBq/LITiikeZu8SMjLajBpl8HSOUIvjLc7IR
avu4wSgmdQ4QB4UGyuLTciag6/fdh+DGLXqUNNUjCMijIo2sVnbQnqMgCpa2/1GfKeZpw7q/MWWw
hKaCcbSFfXltD65yMuOhSZvUfQ8wPPwKF6BsGoZeczZY2QLJXQ3m/nyf0sMllAVc8si7ldWFMBU/
SoKgSLKt3LVFuDsa0R00LkAldqYW0WA1h7tVDCv1Ru6UV8pJPyjmNfEu3DIHd2oO29CwBM8WRS9s
ElevM5kfOr3nzT1otzI5E/j2MUryOVci0nClihSknSPxkdAsV7jOJeylEVPEq8ejKC8aH1W2XB6I
Sif0k4WAAe7ROt+LzxCpWG6AG3W34YA3wIhlNbiKuV4IB0kNvtDMUXFb5IXVXNsDq3BWYUOcqhiZ
GUHf9dhhSJnwvi4wgoinXvZa/7QlAZb1Apnv9VoGobRsTBK0gz4cJuKwM9tnFUcpu4//YhfqMIYK
1AZwIjLNgF82m9k0EdGPD2+LwgDAoPh9mcXYNnWCGd1u5DE0u7mfde5v0poZBwPHFp0LOBRuiw3N
rpqwLSDzMJt+1zco9s1BIkO2YT9TJgz0hjguAyuD89xLoNJGhpEBJqGe14XKIpzDJ+tY3huKHgi4
cSvKkeiYecJE4v1SegSPRsZkm/VXxdfV7yf8z+VFV6jNmmAuS0UEgVbHoV+gJ7clWnzLV/OG2UR9
SrlqUBAqP6cSd7VUbi6WhDCnAZZl1bHcKur8YpaKhbI8x1Aou6kI5qoShlc+IcfDF7TzhdWOALVp
T+F9CLJqWsZsefWhlx0N4aXblog6dAITapkptp5Ro1frDGEsn7mTr4+KfobtRM/ymZ+MYoZ/xbBD
dYxW6335446d6tAAAwRFbJ5+871W4LpO0UFDdkd2iDhHt/35r/2U/ck45EaOYcGOqWroxzyQ72MV
V0nLlAJlabkf3fZFL3VHu/oFLsgIqz4dq7xiKxYpG01dhODx06VIxgK5PTj9Yiw7UWsSZrq7mCZR
I/oYyXaaxdbIvZCwYAFhqjeaD3/Vtrlgi5we9T/WN4+z4iGF7VUjoMmM5ruIvqV0NgtvUK1up/iv
vB6NABPmPLcrUzlOJIfg3JrPNtQU8bG+JoioBT0TuDwjupQ9NHWd2aH/VoytRrlEKwHS3v+FsFIr
l5enE4K6c+Nxoj+vt9aikbXF0PNrJWB7FU0M5gx+0NtVgfC2W31WTAgUuLf9PD7w6c5aa9butVgj
IOOTGPhKT6mEcQYj9aRyGgVLfc5vDFMf9veaSxJc4pRCiJc6FXbaiuc8kACYya6yGzI1cI4gGPCB
yp8ds9cZlh+JbxSRQc1thC7aBbKDpodLkEe8yLOw5iplru0e0ss8Z+8RA10ZZH5crys/GVWknfBA
1i9ybYMWTED3PQ7PbYFA5PYT7Iay2NupeNA1Eq548nQgq+ZnXNQhO5EQvSa9Fitx91NcYL3il/N+
kkbnKj25fTDvWlhLZ6EvzP7Xvcb5O2hAqobTFxFWsNW7u+q2KggEkEai4vcJrixZvj697oHQGREo
KXIBt5tWTm89NPAgpLKwcURjET2z9pKFrLqp6qhGdQD6i5sl7pfweDkGOhb3IMpEzFivSg7q7wM8
+O7MEidzxkgWe7JDZQG6qKGnKtcJQqYQaycKbbLmeBJYu94dldhhG3nTkvyCHk5cZaloH6fI9JjT
HIemrGa3YSH8Q1xIB6kjTLXZNMssK1xHRbfK9S0tbEOhp9w6YqopUFUXovAQLLYLyuDT8ISTKAeG
VKRj6/mAW6dAxE9FLeltD8kS+DLXyakM6Iq4XqKze17OgTfWj+UAnCJYOSqFRgA2wMpgSYjH1eYF
7w83hgFKha/8ACy9qygC6bXwoFrquMpgkoENSn1wMX0fWTPUnrk7aViL9yyxGoEMxdR22gDdgVPl
SnnbK03vomojLms3z/61D8z8EF+O6NMLq2THNZWi3BRaPEwf1vxc48LkMiXeJ6wwiEhPjO6a+kej
5bVblpA6rsy4KDvCdUKb97tfyuMJZo5QtjAgtWRlPecRWBI6u4G/0xvWx/dThfU7aKmNvpnSiJJX
sKeypzZlR3WrRNg9NKX8VTRKrD4YeRqG5zxOHBRFbeYrdVikbme6xSvANWvdYMP2EyL8tpf7Zgdz
4lEQe8lfuXih7uxsNlSwNQe9qgeTLJ6d/TetKhnPBfy0lT/zakFwCx440mlrGM+n0PmtJvsDW3F1
qB5HA0tkEG8PhF1XfrKRhR1K0VFVtyqU4p/Buc7oCdrLqgZsK+2JSJvL6P7t/oAqU/apucTmKwRl
OkS1zQFsD13zFI2qxYq5VRSXe7GL1YPQzH66b1E1ZxA7uSEPcVythDurvjRw8VYhA/U9KL/Kefjy
eX0OfWSiiXDUqauDDaH78L+Fcmfgewe0UGMkoxDCvgbOGeA2rR5M2S5fz8hh9GvoutDY74nWqNzF
L0W1Mt3Aehbzrw6yCQ3JGUq+sU2fmTN0+lNUcqPnMtaRHCYdJzAPgghS5jUe180lPUyJ6khWLS3n
hVbkIyEDeu9xvsrJ0ZgE5lXLE54GM4HlQY+80iImxtL/jcQoRfD3xLDMYpruK9wZbKY5NDeCjkVh
d47hzJ40gOTd3mVeCU03BBNSSy/63dzKDzuTGjWSXHPYLxFTwtG+qNWz87c2xk0TyM7hIgXwwXZJ
casGg5Wy2hfLW1SJrpwswc/SvweFsjQJXHn2ybrtwgFfVts1Vdazs4m6HOrl1eZPVl5ySgIpZetB
FyLAw2wTj2SENspS0k6fnsLhPnOepgxIXpIJHw2yDFxiHbsnpM28NzoFhlpBi8eodqL5P/ghKGJm
aRJOg4S0rqjBx/qOtK/zUUA7Tnef92mHvihc9w36H4YV8SHue1B5d1IfF3U2G/FjvOg3QcM/sAY2
K+UZv7cLnwjnb8Kp+ArPx98+3BTTeYcz8GAmdQDLGpE/rLwsgXO22seCCNmv6P/fnQEmjJh4QrGq
Q7+ZewjvoYlvQ+KLqVArLHNHNMWEjA/2xDBNqhOo3zmlM1m6dNN3y0a335qbmx8ZP2g5lv1qsQul
KEIw7fl3CfS1DYophA6mIsXm8XtUg+L3dg8+tfbko6svF1ap9GuppUTi/HoyB0bB/Noy+ohfQW6O
VQpDRr+81LFFbACdOf7YfGZBGDWLdExyKT/GMerJu507J6MAts1SD0vRyJ48iilIeTXSWh0UNuSX
BkEOG/oxOr+RX+MExNYdvPS56IyrLZ71rLGRYyf+hvjNTA+DKxlS/1cT0xU8zFcxWPWhhTJsjWjo
OUs+FwSLrSLAe+1vLyoLyF/u6fZTX9VqG/YGMjVlHt6BujcjSy6fFBOO5f9hd5fQjkfiSB6biXY8
HDfvge+HtF9grSj8WkK1oTd2BzFeBuQq48/jDzDL0+v2U+fkR53eSn1Rq3TusjhfPB7La/ca3mEn
74oPI3EBNzh5IcemKu9VPpTJTwy3GII0pEWVq3Kkrgd/LELPUR7vPkY16f1boBKeys3n1CkMr182
sMLNGc4lwvFfDKwZXbuVdfzWfkuuCmYWJguE8bdLMOUq4ZQZohZYlq0DXIoGAtFYzRkYw7GNsIFp
MiUFo9GtGMt+Km3sme7Klr20B2MqUUUtXKrMGaE1D9ZckTZc5cK+CxXpA/rnE2bhJl8lD0wHUl1F
xjsQzOYqklxXkjSJDDD9nRG/5F4JHZ66zfPOwX4aifXFUZ8hFaJOXKDCd9QGp6euqR67ziBB6Tf8
4bevH+6KRZfo44TbloS4WqUwU8QAiwPJ9Mcgb/uquokDA2V0tF6xGBuL8NxiJBxRxWYkZrFHcqUi
M62YPKKazlvz7DCW53XuQ1TwpthkmK8qkKUOv3OvxCbd87dFU6Mm1vVbPvIegaizxrQI2dFzBEr6
MWv5mYR3naHUhSMUxPqLP9jFjYElp2YbyMv6gG7P1x38nkyNFC+KTu6QiCeg4SxKdHI9PQO2sWN3
nXtswH6M+EgAlPh499MK6Gdj9LYbPgs6uRGkr04gsuG5O9HmWPTNuQCpJCkN8NPhDc8HPwyfVwC/
9PjOmiKTOAdKqGvxCGUhHCpEFez240TTUWnVrK3Z6ZTVfy6go0kZQc2ZWW+eLhYRAsQLMuwnWZQV
UYF94KOhc/MilI+NZnLb4oKlWYCFxjGU+GCMVDkSh6eSRPfPmfoEY/Nllw16C37iWIRDXlUQpXQC
waVK8ji7XkAKAaxhRHETRNHnvH2gG7Itl+g1AVfKCIhzbDriNrbbp7+IEo9lIMhtb8lTppN6JgLD
k5cc1SHTe85scXdcJoQMheiTPlDFwBFOxlPJvLBxIuvZbHBw1/bpJylmZCVpd46aVZ9HyhJseUex
TO3GOJxpZCsVH0Dgm2dPHMda3ShKtTqJioqrpydA61G+ycrzdjPYtFHmgbweXkSdVNhTPD5wrj1o
LQMxFbkevG4hSRlThdmBqKKZkUuo4K9m6el6zwF1W9Iy70aaZ8iE2BG1qMi+Yq3TQhJIS2AqzNQh
vuUku6T2cThuKVHr6J5WaPpUl/T62ZMWI4W0q64uQAXaUHSL3uPIsybpygYenrrx3BvjbmBO1Miv
cdHnC/NV+5iBzq8+4vC3koH3r0wqc0yyoG1A8NWPoCeVodJQhJzw4Lq599JqE5AyifQ2ttcojif5
Pzq8TkQ4ribgWVJAYgmRlBwMuZJDu2JrUd6M1+YpENxzo4roO/oZ7U8u6aoYyQwHiHGF634D3E/v
ASMNZhXZ357UNEsO1rn/UsIt+ybGUvCHbFYW8wWozYhXEMl3vjWwbAFkHIbkwLXEOYFcwSKd5KsD
d+c6VQrZxI/0+ckAiVyQn9ZmaAkHoztF+lWqfcAy2xfbDGBBgeNgFd27B6kU+CLmp5lUxHR+7YUV
HxTX/BjZehthZrX4BINKrt/FiFmHE3HdjpSiecWtYJRTc4pMeUSjrrTIjZ7jWbopSocg/9+nCByc
ybaplAqWvKKlsn3KbH4DZiJys5e+ltz6ycDYWS5mEy281o0ddBhQ0Ha3GLssyL2h9Cfp6HzLJ+ED
H/5VPOvMYAL86AwbvLC4dhE6tMOkfmAEpzXdwirOsCCbO+sTxhpyiCZj6F10Z9muIty/9IndW8cD
FM3fEK+dXTDtgsFgZZ4i3weBwPrZvE46wPY1iogZFj2/HC3Dij4kcttWjp5mjtaT0D51aRCWN6h0
NLczHi9QQn4f8sVNStKBnU68nMvF7otmWRczuaJcutZwWgzvq7RlXHDgoiQgm3XVJL0xZHfgVHYx
C8X7aHmNSlO8y1y0BYK3ggCgywFbHR8zjMaOJdNI68fwBUdUuP0f+hlgRIHFWhA6jh93My2U1I7G
dn9x/yfSz8pRS088nszoH+EC/0D2FOVKtHUpoTzdkf1mBz2ArLO2Xcur+f5qeDxvnmhNkMFonKzq
eG95DOqtEQJcNIPvQm/thfXt4MvaYpy5trsozMBXaFMZxxyxQE+qqNM/vU8Ta+Qx38MFNa7nvIYM
yfkHN9TD0hkUMsnEPFN+KN+WdWbn8KeMXXRBMMLDLbaAbPcwtk/mVSHZAEFKz2tp0nxo4lDRuGks
nUmKNDGcDnlcvq6nk2GV1Hhvts+Zd0vqM0TWpSXqj0P64g3tWNP0Av42wGNj5u33aJMWnwPYsi79
r3T+wUY5xcHG4dSpGfj3GWzrYVNhlmpQ1BoOdc9JyQ0F2y5qo5MlASpG+Pdn3f8a25BMCliL7vbd
X7G14H5hIY1hxpPaaRlPQzEZ94sc2ePtIfk2XO4XeT0BHMXRl+JtNJ5djhgzTRum/jvMS5UmqCjn
oggLLDO9NR7K2gbvJk4VvLLzYIBqTFQvhQRYcwAxqmlJapT5khuP++GV8iBCIIrVJPuNOPdWt0sr
cuO4yrDcuSKXPBhzac49Jeg1wKaPoz6VDOib36m3swtNG+vAjyHY5zMFYArsycZ2HRpFFnIoSQlw
XffKeSkIw/y8Z/cLu487/D1PkSuEwew5r/JPZgG7IzhsRD7TkAbwHs/aesDI5VQSvJCeoARp8y2i
ncJSd3ZudC5C0h1Ux0MKJ+3S253ImmvWRWJlN2B6JnPoE1/OXGCSGxrm0cExSfoQfwLGaDoRcxYE
HugbOX84AmolN+pDsT8o4CAZmT7S47V1B2UEdFAn1/L8gTeBAI/QmCnsEhmAhLlCJ9DEIOqb0p+A
PBVB7VSwK8JtFLUNJOlpcsmALqn4gNQByQpp9KtKibqKWFPXA3TsnVglEl+I8BhWYrhMU8XgtN2d
tTuR7DWwYQVdR2wdOpc53i2GpGd873GE0vPdnV3QJ3k5HRsuykgA/Y3QYFEV71xMXAm9LMD082xe
2hnAC4ca2NekNo8vYoUQChSnRT05tJtqr5h+5FkTrreF1Uc9USvOWHGOLTGaKkOHep77I3jBEpCB
rxeJj+qJJpGq48oWzq9FMCpJ4FY5VZVkdgIa1PDpzM1Lh/qLz/aXrHsslJBdk+5svLAMR1geGk+Z
l8SqyDvLz6+rQSiZzZQvpdl2i9IpFla7te0LohYrmF9l6tBvxGhjj/bzKQG045BwwRe61k+7W9Gw
AQ/6AGUSuSb3LslfR4IFsEKFhWTBsx+moJH5ce0/H+D29dWCJTsnCkL/j/XMyi+q3WnxMQs+R78n
2vpvvAJgdtTrybV1b7QSPpJWRCjRhsiKP2/T3EVsuedJKN0FM3cmlZCt42LBFaw87nCWDRj8Q2d6
TVQ1M8mN8Sy4pFZ9kyNTN0x1mDDfHf0aMzad6E1IIKIJCTj15jLq99LaeZrmJQGgsSAUqsbnTKGu
qTh25W0Clz5znssT/8N/M214fZcnD5zugzyksudaNf9FErDCgPkEaaVw5V0isuGlEe1d08XWY9YY
WKD+Jfd353m9AkWrrheuwwk1fsofqXWJfRxOEhSD5WKnMLcuBY/yehlqoIZP3MwHNOcvyDegFuV7
GZyZVOQX+YW3oznsM8LaMMASBE7CptZdPU0KjCFFx69Ai8RI6EUp8fFnCMFq2DeiWCCEitmFZp1J
iN2zd6YjsPOBCqejUkBGqjxsjrFwiVohbQ9ZK4L+VJtV/7EIr7LcfRNR+NgOrSBL/i11zh9YqSht
aiVrZDHk789WykSg4G6KYf+zO8juqk4fzgwmowTlV5DUyeiQKGIM+Z5UuyvRreOTanRvs4+aqBWW
w6uvEl6NCUCjs5iXWZxriaA2o3PEgQ3HN4M3GCVKx24xgKH4y95jHH16xMHGZA2Hit7cvAm42J6x
mQ+45ZlFIe3gWi3Ja1rRW64Upx6K38+GvFT+srqHGXYzhetMha50sbH/lSuZ7bmJe3CbgHleDgSt
x7dhR93p8K6SN0CcpofGVLiM/kHgUbS4BDiQ/66C5ffVfBQ1FVYIQbjZZyEQ+OuymPzPq41CfLVf
4tBCrN6rzz8yqIQyIYhl+Zuykw5hKz4OxYWILg2cVKokj6+RHBU6SS+omtBFsOhIeFas6v9OWSvg
ixxZnNGGoS6lODwdbGTlz0rH7YTSvb8hLWNzjwottYxESY/bnkPAizYia5+o3IilBC9mRVmigtbD
kbNA5Am3BlUYj2oV7GWx8z/rLKdvcxg6644y2raSpIwsdwa/6ePf/vSE2UP0n8KNaJvRDpycX+Nf
D/fuwSCPjm1hdAjvvW8IdxwOh4K/rucrkbVOrU3BwHOiBWmIsA3+6NsTRx6Xk5XDJ39LVHChDfZV
JclIfOrVgMxA5NWlz+T5Tm6BpnTSZIgDZdNyozwG7yBlRjHpA7r8zkXo5oZ3dMehrpxVF0Kjd7si
zX5MoG5Na5YAMdFDGfvzAd17oiymovs2/7XSiyjimqG32WCl0LsaxOTGFeJbC38pdr3LHzz0k88E
uu/nTicgv4QdMJYyIo9UCczUBF/Qg1VKU8MhNw1szcA/cCJvP+9wfkY1gOh3Ij8DyHpBfLJHCCsH
JPxym/0VBuSvWcg71If/CNMmFGKZiEtbB3HDo43WLKixi8iDTIW2ZL+VsEjxtBzCqWBID43yGB1a
EaQmGRsLV2DE/gnDgDB+1L4J1YF6Mvemiyn2LRw1v60I9Q7pq8TN+N9TeJJYq/bLO6NWLsJCvlKZ
PeqSYWzzHKvK2H5KpMqlvakVbuFkCOgxn7Wy56J5qQoYENEwgM4K77Icw+P5FjwXH84/z2slhhIn
QXjsqf+75xzXKp/qQco9zj9dp8Zq7UdhQJz26Ki0G/SlgfrPkyi8mQkSagEfSAdBuXw3GDWjVUn4
vvVEDj2VUNflyHsNBikfCl18kE6WInyk5azRrMp006eQ1PCo0M8cc4aaQVUn9c8F/P82AZZ8nqaD
vyNOF6pQhE5+JzGlRFeYQSGzk6aM8ce18kLg34CCLGmIfQr6YAsLonGv0dTjPS26AgLx2sKMBnUk
AI1PGU4ZVOmoFYjnjlZXwSkQAXhzwqvKyolO+3fG6EX9CWayhRHTDdaDlUSAoEChjEc2nlfC6eHK
fWJy2snwE2dkbLNdKwl8vedAf9zamehZMcz2Jy41WFYJrUgzAD8c4ceWZ12u+AaU9jm1g2v/hO5i
TivNQ4UHOtNPypVlRIarUqMMqx1e/0l+mJWA6TnEwMs2AYgb+Pg+/ImK6GNO62hd9wOnvdtUGnQ6
iQAr6/mXLltK0lOHyrIF3PGTR+RY6eb9GD+l7l09njBAIM4ZyLeqyhPh4jvDv2HVbOpLqskOvDkL
VmHnFku4vUlfXv1IL04hzPKDxe0BWgORJtQgEI0FQVhif7WRDFj/tiZP1SqmoCCvmwTXpfLzh8dS
38UTEcjljjotLQuv7S9oX5dvCHJYub5S7QXobnIpIjDL7h7W9GDdKuOBePxn2bIDpXMzocPMlzSW
h82UG7JD5/lYoqioxntpZRTSpAejg/3+OOhwh94VHELcNutl2d9M+/yZ3b428ZhYXd0TJ3+jmLIs
sdCb5cO9VDAc/z6OlRa6gGOQsK9iVNBM5k62SSZk6Nowbrg9WlL/uFaET0FH93JVse8W4kTZs4RV
sj28UCiziRrgDo2DorJHp3FlcnvAP+iKC+xpz2PacHM9eu/5BNn6CI5spsSiiX2KxJL8Txg7Gw3e
C2tReoLlYi559zxY4OXgdtAmFcULTlJGVyTqPfnzRzpPRkJRjbEBmFIoyY5y5cFbaA+1vzjO4XCR
+sgO7eamldTWD3yBoR51s2BlUpwssysCNngZuML8KvxJSv3VCBTsvDEyTjpHfbW0tHxBS+mQOAhV
F9D/p2G4iGQut6QRkQiBzYSwCzX5xOCCOg5xy+TL2xszaxqJrIy8wGB4aIXMf88G8GSvReVzvAPa
RqxJyNWDImggq8dBJaTKkKuR4NcKnCZ94ouW/ZPiQYsw6dPoHdb9vZ+W0WlMhjSI5h8LNAXA1uk2
3p1N9RzSTJqyuVvFDFNq38U7vx8iTZ4+VZS6vv2tQW6Ql/SCvNM6qsEgqhdppwcVpt5z5vreH4Xy
KxVygxGxWYpbGHeOiYYaJSkGTBrV+uPIMxaNTY3etS+y7SHg5r5zNrVuFUzuDzodlQtzfHRlJQxT
lLdsDPLDR69l1DDAmb7zbB1w7l9OT0rdGk8rNEva+cj8qx5OEy2IVGBIQBMU3bw5Akm5ZgE40kRq
5MvXHwW8Q43oWs9NNlB5AkYBwPq95SiCq257yGHL+s2eTnUSOTX35nReTwyxjmRxfLkVVIYuNey2
FK2TWBP/IH88HM0iTz+jiJmoOVDZ0atH8cbRy93+yt+CAr1AHvTOC80cWDe9oSKLUUqwrlYVmHqx
Ec4mOU/+V5RdNztd8Vn8nqWpZW1hr5oBVox1DaEYU7COoHqr/PVtlJFVVPIyoLAQKhe2CaFbljur
xKfaAl6V7rLC13h9vpwVIChpsTnfUu5xqg8GGzmzBBqzSFkCdJJ9fbaHGHJV3ZaSMWjaQeUJjf6j
QXhyRYz2FG+Lth03Y2fZCpdO2k0iZ2tjrS0Sx6s3BGW1mZ4+Atn8evfwAoXz/1vRX5xmaA8V4JsP
RHT6nmOh8NOUdzKhlC/XHwABDrRBaWwtAj10YxkAjRtH/JG9qQyUqozGMBF7cVLe1NnrsJM433Et
kScc6pluVxpRXo4bbt63F8sjfsOrBesYa2XiKpihQt1WeNPMofKR7APzZW+9Nc7TUa5B7q0yYloX
R80m3xMpyKzKt+Fce0C0EAAh1DdBs4jok9DTtHJ/wDsfB/4d0enWmapn+VctbKQdFMrtb8uv/lQQ
NITwJJplvKd9jprYZ/0ci5m95lybH4EgLlHWZAQ/AVP+xIapC+JCmWfqP/aCz0W3t077Dvcq55hF
0hOJwD8ESs+hYZVeqPZ4UStz/qraDxosUCOhEW7HdGL8QpOhkglOAeHA+8rFDkFAlRuufGmechO5
kCWqBbPxK2qP9RIsedwXtb2hsa/yBn2kZIRkcJMTmVr1CdlN1IU7rXgnYz+vZj3ZLC9qOc9MHwgZ
+VjrEbpkB8bejI6eoS1eOx2E38TKLCxH+1URaJg/A1y8BqlS/FFONnrniUwrf/kYFO6PN+Om2xwB
TRx/Ua83Ew2ZKqwVJ8GAemXt4COjw42y8wE8bW+UwD5vuJyqaYuwVP5HN31a+IEmkHo3n5dhB6VF
j6tiggrYXOz2sNJn+GTY+DIdcMoiVyd/I4bsoGwSRV5Yfn/jt0Ll+/JxMWZ+zdbZAhVgrGXrRs19
XV1kWGDY8QfObFvth+HTxn+zinD3CERqsqfVdRwwH6TxITMbrlcAclOCG6YSyd8rBvtUgsGM2oGK
9KOK8xl7qFshtYFTRXVyoctBhb34wHZ8A1zsA6n5uxj0R5ItA9uUjcNDwbEdHWqyF6ktMAzG0FXS
V8Wd8FHwnrnSmw0qpzCALJGbYr0rFoxjTbQoTf3milnb2yfJDWdelg/qK8qJRytaOOn+dudbDNqM
69Rw477jJ+N2U+YWaAgoBFwd0tG5QjXFzSCWvyEYEdmEq5NAznrq4mGRRKntyXDXS5UhUi1e++LC
TTATxQ2/fHNqzttMidOYdB8bK8qK63ZENDrlr9SgcbWZowhWMw9WX7+fFNfd8dgwZMVgKmo/smmz
LRlwGoEoJGbmMV6r/0iyymzvZGcEVEBigzk///RzwxGNCew0HHdOHrJ9bTlqjW5vudngI8jEU23Q
6e2hRJoz5nXFvMW0RGHvTcQwPwUZ08lOSMT918A/7RsouacxBrybdgAIx3eSYZJ6LGvU5v9rQ/uf
8w0jlVuglyfQP/aAvGnyg4Bv8qlLfZksyCeOwIssyvZ8IEHrtUnkbKDpilqDOOYcTViHPhzRs2QJ
iXahgrMX4SCq519hlm++XyA0BDautnAZ24H1S3njM1aGUUb80WFLetp75PAsx4Gf5Pr4vkMMS4+j
hi6DRZ7qBUSAXlpdACG1ZmeEke3W3r60/lpEKSHfgMmqP5wbrTc1w0u4s9NASaauh2VYMQTf/Ocy
yXro68wTExD2gDfMXoowKzsLvMGyLPwAVCyAArDHN8aKMWrwakhf6gXHYCavrPlpyd96RTpslYFh
vF8bh+IW9oSTawvkUKFcTgD2O/2GhOnR+NKt3o+oviO6wwpipbjXseICxCGulpAsgc0feEPqloGJ
zUcKb+1LrFYHbbvEbxJ8aEAPF8/JvsxUUOp54wspYU6k8Y/DxVlCtv2JBMgvof8kxl9kPqoJAwOl
zEC0a8OvI6/rnnxDDGSGh2BgLEHnhvojPFYHHxZR6CHJ6/pqcus/okJ46bkhYom5d7z1mXmeJZkM
AABFUO54EcIq9YSWv9Ws6V+RgmMHgiiqQvPfLa3hQLHiw0pav5LiGOsGaTPGpx+ZrzzPWvfqBW6s
77a+fkz4/7enZZmxHViDr0uZDFbzgST4ugQMxGRb/bOvAgc21wAMEECFCUP1ppoitYFjAVcjG9Hm
NDC0urMPO+eScooiYwRkVX6MeCKapPYjy0VlH+l7nFDacb9jfoG2CDyXyRdLM26Zdq1SNoDi1Mfo
Nab0dAvRDz3gnvv8bAS9A1SsmBJDuJx8sH/yQ3bwHm6d75nQ+G1LHnQjYIEB4l1UeH4vbXCyoQD2
pj+B1lg4OToFLgeixU9RZGlxGmLiAa9+sI86WHoDjEnGpNmg16Ixt+3Pk+NWY3OOpWyFy8embk4j
6uSNpvU07cJ18n0HXWm+FMjpDsr5NiqauLig5rYS+znExzsVCjAlKLK+gPGVivNnQ0wlDJD8ikuP
1Za+3i3Mxqs9LaVUy2d/NLaV9QWE9xxiYv4gK20tkov/bPGUiIasBLFofBIdaER9vskpUE9Je99z
vUjTDTeIJqzzRl/TaufJ+g1/7wqtE3UdguBmqBX8nISBCUhmv018scvVcerqQ4wt1uU2etx0W9WJ
buJjad4dspiYUCwkaLuVAVfOp1Qm+MXR0O6nmrPkB57XTTXiAlfpjYoqdJcKxw7N3LYWoA2rgkAW
66TOPu9l3U+dCVo8/CGZr3yuMORyli9XXsx+KM8amWHtwaeat+NaYTXBJmzF2lUgABpFeJvIUhij
NM/cXh4zaJu1HiCndQIwBjP1r/BjjyHzMw9rUtBzpIlPyd+iJ9WVjLGkqvdSKSfNhceLFznfzwlu
VjoXev4COmCLIRs1F+8jPErs8xxScnjJtfQW3Ea53lEt1i3AY3RPret132Eabflp2ylnwwd3w8jW
UUWi0eUyOfSysR8lu9JVF4GhvEduqVo/H5yjRKY1pr+b2DA10ZG51XwEvbi2xoLIH9mbP4eYKtEG
/z+xdUD0Q5a32CdQUeCRUV4qp8KSl1V81c3aRuyI9/fk9cxZd471zRXv0HuGILWHtFFi/qdz6dpL
fzwYAfuVcmjwbs7caCDb12XVh0ycNqLATxjUQ3yiuQMIRaU06mUdwHQPd1/Liun8jvOr64wcYPTI
ilpPhlSb28+rHuhwkmktZmEvUFnyeGjjfuDC23b43085kSpL27WTgRCkBnsH25OC4kSQ6mnsCV3y
d3HaQ4+ncVDXLjGhzDKPWf60gRSjaPxp2tuZcUIkxu8NSZkVxTPIddcVibbl/BmPMZf34bh6vGMW
xw6Ne59d1mBlzq/e3fkXxRVrkt59cLpUzhKrhtpsjDfcocYAUmZlbCLc8uOmt0goS6j+RMc8DbLV
YO74s88eQZSIgGEfcyZH5XLRdYYGpLEJAVeitw3zYJNVytsLVZXcrhJehJZBnbqS82g3QfTAHApZ
gYXgLXMdz6x+CBrpRykNUsUEe1bghQP1KKRyQXB/wsDgQ6L1I83OM8uwLYvrWkH2xln+hsswxnbb
+X2igN6pXdjB3o8r8krKVSd3pKkGVBgJUya8mE5SF9RB5jEtYTzCu5EGKkk064Z1fSTzXn7gabRQ
UEweT+pGjeByf1OjqyOoBd2itsat4Fj7TUCpB/AVmVQJEtkmKnRcgpxexUmgJwxusv3G7CXyjhdG
uxnuPGLGOmgS/nE8p0I4W8V3lfRm4YyRgpAHEN5XOPdWs+QSD7gWeeNMsuAFXT7XWoSbZtud5V8n
ZqfY7enqT/IbLLx5IrISoTe3dOA9l/t6wVFm8eJphtPQcRC7jEYTO9ZCh3IxltshGQqLFq5ISzyx
JZeR7YgHpf8C2aY//BLPjgrrIoEh54g8bZ38tWpxW29mmWfH5Kco+VJtEut+qShZ0sT0oN6zTdy+
MKYmwu+WB3UhOtzLtNjWRrXsGbjpw6p8ZYqdasr7ZQudcCWFS9qNok9yN1rYRdpi+OVlI5j81ZIZ
Kc1Ftj+WQcM2jKZufBFd/ZjtymI5cNzCTrmCfvVBnU06ErBOrxTrPfAIYAolVMWwbuFYiupkDbj4
qRw+bw7d6Ut4NY+XrisQ/AdSLxKsBTTOQxhWqQFJK0oPBEi/rA35TaYcc4oZ4aL+Sqj9AF4v8sAT
kw/pjHjvmNCn5/vgtZo4p7GidjKDzCqPA3maUn9LM2vQf4+o3MKPVY3/Njcjou6jABhAc3J+gq1g
BFQMH41zs/NsN8gEmPkpGfe6vr7s5gg4Vr3lv6FqrnxbdP0s0cmi5BI33e6k08s5fQ5XpK4p07do
HVCJfYLp6LEc+81h1ii4wHrW62PO92/hGBdS58nLaXAfDyvGXqBDd6wvhCnVeyPlI5Yt1oxKQczT
fvBBLNUg+8Kj6zK8qHcita9BH0xsIB+RO/XMjxLWOpiW3U3wubkDNaVeVpoK361j6wZLqNFB0nMO
H3cGIToTkQIb5EjfsK4fCBJ/HQYUusKRoOo81FHKrvel62K5KwbiKSaFoIKnzljannjonw2f/Gwf
zoZ04q6wcaY2Z1ZSd0SeYocA3DU3czmSAfhNn3p2CpeEx/aXF5qqWeU8kGPHKwnBwMoBY+HjOUeY
Qs5dVWa4dzxoTJRNn7tu6i4w0GIZoEajTDNqGcOeHXunB9C/xYjq+O9Iy1sivf1jInFF8Le2IKaJ
f2X3NwjrbOAz9i+d9SnIr/yKF6XYy1h6hJNj+bK0GiU0cOrNUXLHOh87o0T5nZ3fwwmtcAttfxFP
l0Pli7gsgVFhXFtGMWGeJ0fiNl7hfxw9QxvnPVm/nSTQqsoK3yKK7JB7Kn9N7sT1a0OQxpO0Tacb
9GyMWjIGznUrcod/7gqUc3L0KoGns/EO0U/M/dgJyTIx9sN3KsP/kG9vs1L9FmFjtrSAgD6X4rOs
3LOFuvXRtmAN1xjdRrECNdYkduMXExT3cDG318TqWOBdkUGu1fZxZn4SDeQg2Yim9a60eiPW68os
IEwxliPWs/R84aQogbpwWap86288eQ17k7RR1WGjP04yBUbb2Ry+A/Pnl413cbMFvzZ2fATAJqSs
PEOVk8TqLkCGhuzJE7rkb6nQi+Qux1crBD5RiDJO+DF0touOGHc9LA66OhAzrJ2l0q+Ya1RjBjCV
Jeykqa85sxdnEbyVXAko5m+2aRlSeTEKSqADkOMP0iMAobsH84vQhgUWMu4ANJL3kokfvjRyPP1q
pk4LYZoo59/B7S7ExRHZVpGcaVR98QA93lNZxHGZXzOgfFC2uG4NQQGwuFtAumT0OoQ8Kz27C5yc
SYId17pgUYhhJv2cxMuEolGTBXsB80rrM+oSLw8gLe/iZztmpPNyvHOfzHBpH5IacWOhBsh3b5Sx
5ApwzY2022lhxT70B4cVlrN0TOgaqMv7FMIlhKOGIqwNj50OGsf9FJXoKyNoir/z1awYdNDdr8xD
ztVE8z1TjoCN8hfg/AJiHPcFUucIyo3ttwKArMMSQmv7GHNoacsUePhppfI1d1VIV+nqIRSm+wh3
1d6RBf+uqzaKmCgoNMJhyQD7uZjJ5X4mdz5FNNf8YT6FsSB9FY9yFuzepOedIXSFNIGeoxkVa1Ed
0DGEyVvLHcg7HGGgP2P0bJ3Ydxa408GCd14Ib12X58X9NxJn/egukm1jBkyApkGzPfwjSDaRQyqy
6zHSmmixgUFrzYE9zfGuryP12AuTtAnaKA3y+mrxhZg8pM55UlIFnJlL+rLiiSLuKViGAWcRmVND
DKU3apnRlxvN+c34BcLX45XBpk2UXpruGvg786zp7TSF7KT3FQd4rXHVy8PObVYmLzGsARk/ieaw
Szm/smgkhSajlXCMyCBxleWtHU9ytRbhQK9qk+f1xYTeg7lE0AU5B/FrNXkhEIpFs5t88VQNy7ck
RoqQmXtJm5YwAIemNXiQnkNy4I8us/K1auBL5YdBbYgBYiOQyy+tyXkoAPS3uPclKT3BDnKmH6hi
d236UrRPWCpBn3DXsWjlhLvzofGT5uOMZvGfiyGRGTujpao3OdiQlbN69qv7jd9QmA9f1JP0/A/d
snI4qxPsZSN39rs/OTtCQTkV1mVNBlTZpUx5uh2HhK9NxRQ9VpgjlZOG3JRmcV32A6yg6+Bj0uO6
gJA4Hu8aDS6oC+RkbOZlXIdiGye0HA50IsnO77YJP35shW0q3+m+1qKO6NNh3IQq7ytvL89+X0Zf
tZd8Bo9dQ5IrK/BK6b5Imom6Fbf8N1FuotoZZJ5J1vZ8E4itK8jEYkTHz9nObLMVv87js+7SNGc8
qKTI6KgB31rRGMVsI1Dzoa8v4fBXj+NzMZBtsAfI1Pzl28rm8kOAvW0tmaWp2GU5cHj//z9qEVEi
BjMf0zll+CeAaZhLoSoLDSCRRBDiIux/6gFVDLyXKeJp2k4RyFxX+ftSn5H5WGEi27W9pZJxlZnN
3EWIDhIxw7kOyfR7RMJuRsHmfTOrHS1hHR/0pZhGXNJIP1QYBEZUFVhDz8BY/grqjDP//Af/iNam
tLYyT7EH2zMX+0ins4udeskGH61guhdsbnBDZe+RcOqcIDrvkxViHvN1ZY1bGX/MmLjMDKOL4IkJ
1N/JC0J4MCXw/HJI1zZ84DY5uHc0H9CxN+OzvyHM7hyxdVYwU84Y8JQsT+l+Ptyzh0Uud7EYWf12
tJ7rM3Y+HSgtyLCv6an3vgstUbxupnqKzS44Dx34+HCMYzZRB0pdsQB2KSHLvPuncy82Ie4DK2Qw
O3lraCwq2K/an+Mz4I2IlynSMpHHzT0XsXkkEqd4zHvGp+DxNZHEh/YoQml/3M/BNjqVIQ7+s0hw
YCl/krFlpJP4lSmrw82L1xk9LqdQ5xiMeCEqdWTXMGO2IZlf/6yvuWMrmn2vmJKnEbEtx/3biyJh
JtateEsm87dTJAH/cXbc3EpQBsQmM8YeT83WTxg/dkxR+BSL62BnoZoJNsUkmTXopcYgZvwiPEEW
QfZE9zmeEdjJ1rxqANnsEGhPpgyabTRRrhiwsQyfW4akiqIoOzt/eB6+y4Zqz5BdGZmGOrb99R/a
lRxkC4YQVSf20/brCNjJcrQsewMnT9x+A7AkdnTrf03dIFb3x35FQmfL2hX+w+4QZgGJj9Hvazk7
iwGajH6Nr64oU1xO0VBmBegi+ZO0XquouI1nlJxYPbECOZklCz2fjyjbIdbcufAINXHGMu2jA5n0
Ztcy7IoRV2eondX5ZvZ5b6DgXGsehHcCqjYM47e8NKtAont8trCdPxj+d/1iuGQ14LLTng02+lSx
/Xq02UXMDZI6uD2C1i8E4XAQSOrbVQOdBSSOWQjqmVORXtKjlmsOYOWJDQDPs0jx4zSL+PCka8I6
AYtNEB5NptbnzdBOJAnM/e3ssh7vvy/WlAkwEOPSHLhuiTaH6EXu/Ao63pU31MXF1XrYkEgl5d8h
IJVG0OMBX/Uw0QFdYvyd2UATy7SBqcVA2ggOxmSjOni9daKwUifpl0DDCLZVQuDc3ZKONJBcJqpI
19Ej3+3LFsNrQCx5IjKahavqb4HIpaIWf5YGvuaDmFHOW5cRu0nBqXRCi6fl/wjiteehOBBgzhKF
cNcIrybfLQJZYL83iVb6KeXh8CTwm+C69ne5qtB5QtZ+OIETajVk77BI3I5Oy/y2CkWEQoWSRFNM
stwsVQcTdH3SgUjzBvJlk+v12sIZEXAL99xgSB2DHieStESklNqmKEm/o1ko/5KoGdyDnv50C6lR
TyMITmvrZS4IrbXfGSwPAg/qcSWmam0dv8Gl37qJMkhyjLmlt3VpnttAC2UthwIumd/ucXY/GjWb
GLEcviIxGJasru98uIndtnhCr4wsfLZphn2G7Y0LJByzu5sfJIbqTB7/Q4HlrYIvTnRhaUDFV+ak
tvgjwgW2drtUHPBk1/e14I9/+iozTVft2x+/DtKhljgm4GJNrl1DnkLLnk/cAxdQN0SpZ2rccqf7
yGzk2OT16V1txj3Spi58JYnk2Lcj+wHp0oyakNmOF07qx9jSqeN7jsE1qHZD4UavDVQ7Sp+0urGo
x8voBhRNK7yZpUB/xgtIpDSScRCZsNybvc80HZhtQl3ntJZJpwKgU6qzDqznuUQBpU0nXY3HjuSg
l+cU3G44fI61Xk3YdMpxUEJbisxfVRLyPgae7L8nvJk4PlOjEyJSRzpnt5gWNuDrBLgGLVofFj4f
NQfCkH0gQvpgnCoNiwqd93AMkgq/m/LZjSUE/tMCRNVGzadBnpanBxuMZuUtb/NwwPe2Wy+Ty+zo
vTJzKWCsM5jqs3J3KkmnH+yEQE74OZGcUDPH7HjJxvqmbRdbBmkc7SXKryDAOHq5BFvloN4CxJlK
///ubPZ570mPi8joJtHcocyyuWN0c9LdbRlYeSLmRg4b4ricFYbJVEsoKjb9se8tyrHtX7oKcCZ+
9IM8fE7TdXYisHLU6g9avCTBKSb50egRnjGLnwaGlTRke7soyrhsZCOR9dWQJe9AyjloBbT21Slq
wSUkIuxN1i1zUt4qWLSkbjMzlOYLjTBsjwaOBUgQLriIT6GqRIvOrz35KD0I0pI9CcSXRbgfIPg3
uQJFi+L3SVobhzb/r6UYX1gcnqcStdVAWiHd86EAp1/Wmg7RPwuC1dS1NJXqksKU7A79TcnpKG+k
yz9zwVbArp3BVk9DM7dqFtJ6NpQTerMUkDkGDs3eRCVAUiSLlswjAeC8jfRGaQcK5czD8aMcNcZ1
xSnrpYGYJ2+yanNjJRo/IOa+fnD9IrK0FDRO3il0+ow+t07LYK9l7LQigijGpECL9s8w6+9foGGq
dpabelrrMwpdGYScP4ox+nQkI5xha0FvlOPf2Iy91XqNhhcLeUT/dKSfexJhjKP5UySMyLiUTZXm
yMijwm+4uhxWtDiWiVEW2A0fqujGqUgyeBjZrw2WbsATK+68Wp0LpHZmNtA4B4g4vgrFDMlb0QKp
f2mrKfTXqMDX66evZjExAAZ88iVoHKwvKV0pb0OGBlvB6IMDVR1/uHjZvRTgRq2T19TbedaVgtJr
BmaWHuD7fC4eBWw6BW89ecIqVLuXxiEaSADOnhlvLS6Gr7K8ibDIWeKmAs1jqM1N9djwm4EXWS9U
YH5i55QeTWCtJOo+Y6EPh9mYd0kLykjUQwyczY69KsWAMZfAZPO0BGK1BxRF+MSqq5gBbvv0oemK
QyjI0bysrxtuBmaTls+OFKPWlp0oSAWdzTpj/aPBnLu1OaIkJK70SJ+y67G1CFmStbi5jl02g9rq
95xNAwpS/BS1afINCKw5BXZKiUpao1NjQIC6OH7Il1jTvku5ZMkUosyeJlMsHvdK9vnjdtf602m9
e75GxCe+l/E/0KMw7IkUnPZ2vY81m16hKEuLHNFQ4s4Fdwu6QfVehLCRUDlcrj6LLKPlEo8920MC
ZLUeQQOsteHDHyaTmY60REswYsa+XFCTlSZwZHap38rf+tBuvmXizIB2wKvnVpwUfzjMayyyUz6N
WkGsNJKO9yVgYKAMTRtfd63Jfut4AId17jWrRb139g9ngzrPcCWPxNnog3a3Xe4JNUwyz71xZN8l
buWAt8LSXb3VC0pHg28CUTTKkJriH0GlPiHjcZZQS3+kU683hjxAaSyzyo5xPH5nXkWTUJyqWDr7
7pvzVdJrE8I3JnpsJgwWTSn23Cs04V/2mVQ+d9E0C0DbjiL2VTLBBWxWNUksN5VEhywP2A7cTS6l
TrbpRw3xoC6yyehZCcW3B7TBTeQ2qvjfSP0VNxbAkdnEhfTmlPAsXndvQL/qe2Q6QT4Qwvxuloml
5cEf5/k70F2zjmA7myj3K1Ei+XdQWFkDk8u0g96uYp9GqCqHgKFTwVWiknQVGXL8PxuxuvcviFdY
wwYmiNt+4JFjQn4PFDoF2yVfXXGq5TJoA3D5xz/eSTBG8jId76HNxWLKANjdpyKVH7YjdUertiUL
KM+35QJR2naS21SB4LDabjkK5OMXnfLZIves6EWuWDG/X4GziZ+GkGvL7d3BOljlPvYkN/QY6UPr
t/vNxqxYQOjw/EZ3yyLr0PC9FYk2FUv3B7umfxCLv0GPNNLzHwkAR2Qr40m0VY+AlYPTf0TAr3c7
Hh4iguIvX6rPxbV7IXEkFJ5AxdEOgAOW/PzVmQy381eblIXDZpsh8AHSjudladZ3sHoWdvlEcDNo
fZnezRStJ5uOMc/Sy9NtlJuViJ3h9vn0LJE8S90CwzcKOj6wmx0a9aYbB/1TPVi/FKC4P0QVIaoi
lYOspRW2R4SBlA2zGBoJix40Ol6Q62h0o4mVNb/KL3PHU3PXZr+Vq2kSvKBPTH0Kw2FbnM53X2IJ
jyfnx5hazigL5HaQaJyv+cIEWaoVzw0fkjjjGHAwZCPzrcWqR6H2ViNk6u/ii4Fod8TCHuEfEIII
4glbcmk7C/WOnf4aeh+x2zIbKVBpLswnvl+elgk+m914rihEw6uej/M8DVJZCsckWseB2aqqcfCT
I8nGtCMpvvvuDr2qBwV+t6Ugun8t8CO76VUeHymekTmnvLVvBKoLlnsVVmLf3+E+9mX2Ui98urBW
rRo2uZLxo3pZ7IqsDUC4bMWYOugsswbJ/WHwBxOPv3TwHWp+lxvUCWdCPsiuWBOds9lilCTi+CLG
bXdXS4scFsyqxXBBlreAj5nRX52PIjSjJdlVxP0cuvpGY9t1ftQ9EMqrDniche9DH+3q12K8JcbI
BccnHYQsHeUtDbILOg6U2XRinqxqjnMicuV8qHpEeZ3ajx7A6m1hzVlGlHRXyCio8t0E2eyOVA0o
9Uel6s3puh6j4Jwto0uyIF2EoVAwD1gCNx5HceYwPxnXHQ1PBtdZJ/Pt4mTHQb7UPjXTx/6z02CE
V3ltyFD++OVFmH7seLLVCZUYxm7UZKO0s9Zc/ocmin72KLJGhoUHXSXCIh+f45UMBIoRbIIXjjhp
2NGy7yLRRI1WDgDbp71M7aW1SxK/KdPT2C0CHprLndq4oRUUcR+Ed1tgev1Z8I5OYEmDMf84qAPQ
Xrpzlhf8YLNDMr5AtSch62BfffBF1yRoIDyKmwl12GjTPNd1KDm1Zuz69SOEpH2lUJpwAlnqz4sc
EbNndWsWeWlp5+Otz8x4DvIckK11r6kyfrobaavfiguNGO72zaK9HplMBub/nt+ae5TUAoCCzDDV
yPiPX/osXZqPAa8kDXCRGlJLe9TtupUuxQSX5QbEUWy0K0KS81J8TcLK/ltCYWlOiXsuVY5Ob9he
XOVZ7NdI3Rmd/l3CRvbZL3Sv1eazdeP6UWNPlNMYDIgk/hT6PYBfsuu4YRPiBfYXFaz/cMPEKI4S
U+1tCtsU4dy3p5tLcUuIC9TjT9VZsJF+UAEeWaDIwEyasbiNXu1vt207rZ2A01gQb/4mvrW2gK4P
OFPrMsH4jBMQ5lzrdzYdUwGwtJtSFEBJIIKwKYLdzBZZnhMssw62XXoeMxs3fh0TzgPi3dmSfalV
5YPf/QUM/gcsHM0hKpTCh6Z0Oxo5JWq9RbyqdLGDNycruHpuadW4gA+B2zGE25xv/OT7SkPVPga5
gEAHomYW7474wqqrw6ZQSS4YfBZnI2FKx4e0boMC2YfNY510gXG0m2xXsR/McQ1jq8IFHxZFipwu
9jGTIADlrwgFChxfA3GTAx8weUX+kKDRQ2YqqlDMWrRE/ICFMvsY1CZdN5EfN1qdSM9dKRt5CY3F
vX3+HZpkprql19t6w0IRZIeCflsKRH3WtPpo2I/lWRcoJ9Vu21yDRntftKePNDbMuo81kXW7X+7Q
6qN6k0miLwjGqLWbLUqllHYUFRk8DLlHfWGVvHqtAULaMSXppOyl10FS0K6909OPlWD2oCzvvosj
+0kbB5BXoTmoLFDcZcUOnTwjqI6IVmJGU+beMckmIk6mopFjRLG7WKXJW/HNKfhiltG988xSHhVx
x6/1R/ddH+mFVArHlNwZeIc64EppmdtmXAuaXlbJeJXnh4L1ajrQYnUJ7zqw4aA3OPQyV4slIwvQ
0n3lx73kZVOK+K5RFTd8+j3GX7XSGcBuhSDXveBlQvZlGancLATiScMMvcdLLWQFxns32cCQtsvR
YKNxq0r1G7bBRXXtOdcyvBUQq/ucZlbsFqMxAKgpRci3OdEo87+DGNRV3MbVEf431wMRjIAR/WAz
ohWFz1PrkZhfRGdtnbB3XgNOUjHEydZyx7K40V2ZtkauMSnAYU98KQGaaWYN+avkKREVXoQuvBnm
sOkMxLd0miXnhCxugd1O7eyf/4AtScZk78V0Nm3FT1J567dC1Mt30aflj2xmsz38zqlV3HP1rDBe
odiUPKheRVr14B0RnUZmb/2JZ1BhdNtcCAlgpnMvFF7p76lmtau1pBP9qv8Cyawz4Nqjy+037Y7E
uuyKfYmC5SyMwJ+qtuh5symmJ5zibveYr8BnjsMC3jwS2q0GUpkNrV3sScZdT6sCbtjBa5Mk3oAJ
wkZ8EiDDWJKHLxYRXZm130AhTCmyf3qe5o0m3qpEHOIJhtOey+hV/CDIXqw7U/hfDpxNnklEpkln
dhmYpX3fYlqVJ9eUcT822BYajbGmluClXIyfCw4nwlEgS3HyoHPHK43vJdJbQggGLveNEq0afbjn
LDsOjX4Bl4DXRDGgJNJoesQ6MKudzNJ3N1EcCeerTVe3G5wCLPrqqkRDmxdfnN7v+6ZtcFLk5Flf
QWcgUmQa9biCizili2xJYXK9aebZWjuhZZv/4PpKg+0uOr5CNDHvjJQPI+hY5cqJ653mRf8THG8d
ANcSbXT+vb3z5IpUWMJvTYxs1TuKJ6MhcsD0chpc/1r8SohyfKpZt+I4sqoTrb0IElm68Vbvxjvi
ExtHyiNi68ioGkzF+rtqYtcWNayCQzOWMy2u41AKoPlgHNDf4KLw7mKei9hEtpa6KB3JSj+3BRlU
JrT2X859TXoO8QjGdKI+mPaOlqNdyhqRBNCaM7Osz/xe1uaJQiw9fxJI8IAwYMzQx8ZsmktjyntQ
z9wst9i65S0aGmHFenV5z2J+GEFpNDSJnOV5R6ferD/tTxqbT3HMP3fJBKvWicYay58QZwFMU22m
04W54emHX52iuBMvWrlV6f1wW4cZUIQOMl+oFzikdNga4LIRwjkErTjVSuN4zBWkX+h3dFOsG4Vo
QThcwYkI3Zhsnui5P5xCgpfz1+e5Cdzn+hTriQynj4wyFZF8+/VKRhJBoVMXdGZ44f4v4TDOP4L3
/VW0+zqYIcyTZNCbyNIm1Vp8HXT6cL1psOqfp+tkW5G3YfiIKo/VVviw8axnES3BC+AAkFRiGYI3
JlA4RUV7Tat+cniM265BPvB26546Ms3IkDfziBq6pzJn/fPMBKfx4AKre7z5JA3cSkLGEq60tggU
6JNqBwWsBwbfT+/ZKOGU4t0Fu/9gOkANkK0QzAzT8OJWrBRTEZBOVOoj4cCZw7mVZ/MI9twyBhKd
TuvO4LL7McaI4zS5zrepPrx/Z6X6GLNAHOrEeo55pmJJtF8xBFXtTY29hni8DjTZ+2w0RKMRau2s
139tvjKuXTnuhZIfhRCAHz+FeSAy+2nJxW7gwHuGvBruV0mDcBfs0hQpIPxSx4zQLnbN5yCeIGwH
8bZgy+hqrr/6FnJmG23jR4ObJ/GsYXLstSyTUo/u+lChZJEYJBi1lrmcOvzYEZTSr36hS7Jzk1n9
XazvuLwfG0EuuekBv3gU0MtnIei8scUbKu//DWQ3jfbcwUP//JUHOhpHe1UZh9rzEzIV/a+59oIe
+B7zWyEXztnTCteR/boW5JNrgHMs0BMImf8G+2i/YZCHzzValKBD8sjwfDouYIGxesVgtz9H4BAE
OcOHHMouzyzcm4VvWQzGIPuww9rUDa3xRizyyCQ8MroIDFx3S7wxCSoZoiGio2Ac81nNYN7WaGQo
+8WGEJgtqeab2Ph7UytFL38rwWf4U93zZFZFyL4GABBiLyHYoMRGQsvBDa5HxSYrxLJ3k9qImRy4
stU4KTnUv6Ba/uktRziel2pFgZDSbpPq1Tc1sVEbgau9YVo0f+sj9rYjsqhKBXvQCDpk1wItnjAM
gVyAkjAOR1j6TLJdeJb6js0KIocbuUU5wfd1ajw8TMjz6P3v8yLkemV1QWD2clc8XBe/Ums84QQw
RtEhJQMAndRvxfSL57pEzkPuikepExmto9wbHCEmnc+yIhKae8ycJKMB11+P+Fm7QGn9BMHNPfvs
iLwxERQLSBkSHPoXqZspSAep2os5e4Kp+XMIBgZhDGc9ZpUfeH6GK7NurNEQncSXQFx+DDjqAINY
ZjWw9JRbT3wh8jYhmHHiF1h7aW4xMD+ur46+XPNmvOgW8LWbko+qHQUPCabgz5GfRWDtWNOnn0rD
vE8I3bmc1Fr+PhSNw2TL1vU2jP1JUi/fFfH2xPupbv7h7QO27Jtw7I6dFY8q0QX71q4L95O8mmrP
WuI14hgpSaxIVJIQ6VddRcCh1sZKhcz5A2tbY58oLDSt17decpRDz7QR4BXngz6njFW4j0MnBgvZ
EeNhySYPPnh7VgfC5jjztuEXulM05DEBjpfzcwo4Xj7wSEooiyAV7D+ga1ybCudHIpS9jZvoI2W+
u6FQVFYtSjkC2vvIxlEpIz6aIYgBsImpUelpcFKTGIGdAc3Tk427CVWD9lSyITzW2E7JhnSdGYIF
rveqp2FKOqkMydu4LZeBVecNjvO0EUKuX+I34gYMY8YlD//cuAdRvgxPEQL8HaLmbNZLQdkT3GUJ
1/EY78JT5VAXFtR5YtnA/tItVIXt2g+qT57EXFm4SJNhYOSyMu+jWJ94dfmVKLJgfn8M0CTGMlhn
6GqSWd1DMcPG/i2UkBMSM0a7FQ5Juft2Q40ILjCz/W1SQn5VHwn+lVYfYyATc9+Qvn85y5FCesGB
mp2PM9IxImUOC80gdGVcMENYz/n55FU0sx4I3xb8Kxspx6176g4yf5EHuBqvhlqfEr8y5UG7Ys7K
yBjDK8wjxX4KHddLchzpylrOsz4ZnKZ7DdgwbsFygDjqAJhpqVqaMnaYI12DK5tDCJjafzGSW7/f
15BQV/BUeuP/lzQceNCnYcqzkewwOTD6UYHudNva+2/en61bhW6OqFfFvtlL0/4QeK6qN2cTdr/p
cFG85O8u3xl3Q/70tnSXyWCT386cAJlJO/XaatxXgAqgg6Um59U8uxWL9fVLZsF8rkmg7qQaeiQb
G7h2Uyr9/+wNwHA7noTSUPXtqpSVn2EKN6q7AD30LJAPvhLVZkrXlLb6It/Smt0mVSAxBP0ilmca
AVM3xkRx16RKbfe/6xdvhu80V/A9dYmmY46iZGf4IRo9TSXM7av0V67KTKRWsOH9b9P+4Lo6VUbp
RI5FEKXwzdvRy7NXzYUNMQG6JPlwwJMn2HWHEWk4747glKyUtxNOtx1+xKMUHHP15GbbIlQOKSTW
NxUrYWEkA+xZRSg7dSrbfGTQfK8jwkRou2edOmgQwdxHOwqtdm7wwYze2Um/sUh9JwZOk2+vZjKf
EeW0Vvmqk5eWb4ysr1722CICUBP2zwYHYmF/18R1HMwtzRlawaxrilTqb0+6SqIuDkCvJEhZnhBQ
GlVwKJsbesZGH+t1Kcvhk3UNFhprCR+xyGbYygV07v6V7Ln2E3tHPfzZKMjM4GKD816u2/fVw26H
Cm0/jwrrirnNxEt/d3icZja6V2pzygEsPqoo/cdj0UTH48nUYP5sHUUlyCZ0NGxHDp7/ZhSzK3LC
GCxiceE0TRqydS+UV3OON1twTMjBkh5SqUTxlUQYvpxPH9gENqmVHGvPLNXpvMtLUG3wiAS5cNTZ
ikzm2SV0WwgZNAvj5PoHeUM5RJYxJ6uEuQDp0NIIJXzU3EfmytAlPHgQu1qgdiHQdxBTEsOL6r+Z
dAEdxDKFot92kug0xmE6fxyZl7IadIss7032mzfSEboiRcsqph0xrN2yGcSizpPECkz3G0I4kLGr
RJeZ485KgCMUDNDHGHTdgn2Uki+dHth0EjPwTFjx+HLjxrU7HfB8RGi3daT/Djw2GCMb9hxNMJ0o
dBBoCffVBbqlfrryZVtBO9Qv/kRSd26VLhynFpUfupE8wn0D/ZetJX4LR3FLEPBqHBKUqEREs3b2
D+nrOPAk1uCVk4yA1Y1D722UtAQGwJ/ItcJ8j+ckD9NM4s5mpnaZheSFXfIA1YLu9mhgUk0BaCRg
Uyf5KJzw0rYVggfKwiM8VoH0n7K+xtFdaVqi+o+xdLKISgfl+D5XFpq8vFl+TKrs6jWiRY3ghc5J
oZkjIxWRh9Wu3WSjOsgYHRd7eye88lHhwK4bCmkICFmXlBtY0uGzAv6Ay5vPN1rYGZvFmOmyMalK
NqnUk/kgmvtGnJFZ5NHAYdgPBNipqrT9ga2hKNkG/DRhhchnKGQhW/BpbDHx5qteXfOjJwv3J+Wj
VtJ0XLat9ysQck0qvKzBVuTftNYSCZN832e9jUsQqXRdvaOEMutWuHUSNGPrdOw5hhxxsDoBZL+f
rEGI70tTpAwLmmMo4+BNg1plxAGkEuPvxg722EwFZSXFNVxAhnaRzY+CsiKngzDlgUdWPaUDtMSA
kyBsHDELDs60rwhGnzhs7ztHlNqpHGo7nvLm6HixH87TQRbg2QSvd+gJXCMoJsS3hLuzdhJQNY0P
MW/qnL3X5orN0WP/VKOo9MshByCjAHI1ipDH7KeyQtkgpif6ts25RZEalRbNUb5EPp+8kw2kDWOm
pe0EH/hViXJ3H1bg8eE3DBtuUA2wMGsd11NlI0+bHYfYDdY6wOHH6Ek4T0R/RMuQsMYwz8A5d1dz
EAdNhw3S6xpN1CzujGpsfZBpLp3tI5wv6kJ0GtitjriLf/eyF5FYNx6o8EY/Y4ZcIBGclnCKEyEz
G7vy7KgzA2OTOcW8B3qaWiIJhkFXoIg7Q95mRHeF7ff1i6X6SiWESMwe71427vMc7E6k66hfw99z
lnJBX0GdoRm/RUbjC/oIyvbpx/S9OTvXZ6x7+iY6NGBMmElett3XtxjXaEU+/MVaFHvbh2r/DNOB
MqR3mrTdT8hXr/ug+4QLecbngXcQW3oS9iMeEJDdPzCnaNw17wGxQOEPNK17/FXo3BRz4bsAjIRo
gJ649Uj5KXZZotrZxZVBU0W6QAtLVae8XcujuOnLHwIb5Hj9ew072wQLOB8nMQl1P1tv8utIjtUA
YAB+wuUWIy2IZROYTkV5Wq92/CZz6LF8+AizrPIaTcWbr4WbFuCAVflnyROIZqYCOvDGHz+8pTjB
hbdGfwcrDgmmye8OyBiTqu2mE7RHxx+rijjJNhrpv8E3f+EzR9Sl82WclWRDJ4Ba2X2+BXjV5Fsc
VgR2v7u80jaYPJFZvJNVLT/aNDfTcMSyMI0fN6GrDvy3MyeoYNcUm7/NSHGZOI1aK/Q8SYTVpkZD
1OL0PqMccH4q4AAIhOVnMb7dyJqlg/NGdFdO6iv1mI6qdnnG2q5qgt2HiM3AI/6vw+svHsfyy/2x
Q9glG+nuj8Rc6rGCyXmOimWv22WAvLwyWtdxM3OCL5Rv83mcoDguRKhw1sXyfMcw6b6V89vfm1vI
0SxjP3iqp6kfIFZzDoaEjKTCksdRx5hgdLWGgc5WC5oe7OQwtXM3iRM+dC5r4EHYfOZm7zDCZXc4
R97ACQFFn8bzbhpXNFIjcbCBf/7kI+BFWxi5v5OiCVG5s78BCusHcjIjnMTQYyApl+KArSLkSOYt
yZArBJUfZ8Pb1WcMtlILVrr6x1Ld77P1sZpTSXLQzlpAXAb65ZiuRpbozFXFLgHopcgpkMmx3fd+
goCmvShvLKRp/4RcXhvqJhgX+8kf6N0sfQjbNkFqb4plbKDvn/UHDdQxNBEFQY/glzGlcJLyV2KY
LlNPjgl76jNCnAzmUqktWjylEcK0XBWb4krL5935p/C1poiL+xL9Z6UerO+cAfrYKFR9ScDCkBEM
Tks/WB5sQc4SBlE+VH+4RH+GvNyku7uhChHO/HeOSUYEAOT5e/b7R+XMvWvQW5sEGRgKYjVWcZqp
zb25pp7isypVd8Rl1yHHlnDYWvnk+r5VaeEgucaT87aSk01XNNqRuUxanbkpJG4AGYk/PBw3uq+r
6YHM30x2/tl78Pi/8HIhz6JogFCKM5fsGD8vRtbapfqfC3ZOyHRsfh1I9HYUxrOe6ip94IiKo26k
juivI4MBIHt1705OQo7FMMRerdV14MinUeZt2eaSsT9G1qXIpxdJkx4HyU0wfjR0F35nyjVx+S3t
B73vNKOTBKDO2ulDmtXxNx2UQtFyCcMaUffSBaWa2vSh8ZaVJWCkpp4vOsMZJFIMBoie1D5eWJR9
4ZZakV+clSftR5bmHewuS8p2KIZnZvzBzK698r/jbJBYI85vkg8m9nR1lkDrYmKuJpBx0q++zs4h
LD3g1sOwUvXMtjGptYts5x5KcWkqyv2TVXINWlmiKsWl3O76XI3J981aHwZF3wbEP16TLGUkAuBc
fADPdhdyv4dZn9sRZ3M12bUXY55DTSLPRzCskFRplcOhpFHnC6Cfj3pWtkL0L2eSuDr0tYsBVC3A
q/vEZ+TwKlz4nTHMbCpzLrbQCDfzQwL8LUieMrTGz4HwW4+mRoh5zpyuRMym3nxyV/1N2scIexY0
pFRKqwAvcpnDWIH867rg+QULaJsFMH6+HIhKYFTwMgqrKcMVcN8Bg/eiosSchdrq30NN1Sm489od
J+chZRZ+tao4DOn4AgUGTEHwnZYPuRMtqzmH5t0QHtd13RnY/UgtbznfrxmE8SbXaW1Nh+Lpc924
I562LI310EeMyNRXYjrWrbKV2B68Pbz1C7zyPD9/Pm1g63h/0aHTUELVwZXMAVZ9QmDRjcIgLJHG
wGt2xmrsbl6kDuMEApcl82pUgej8vq5/M5AoCROwPjLK8/t83VmhMrRrErvNRhfn04+frsAo0GOz
V9qRHE5N7f7k3ozQRTDrOfLUb6UILM9L/KrnhnifUkait3Ct3QV0Z2O8hhJ8MPXmvuN0vgSRe5DV
u4MOo3PQoMjHTCxTfsJulr6dc1qSKiMIVYQ3/W1l94YF6VGkQn1LVoOUr1zfGYCwAamJMrYUTbK0
lY2/bbNReNt39Wg8iL5+ZKJOJK5gDTNaK6kF6alPkZCTLTaZXpNyXlZXN4vLFt/x3J7yKdA2ispH
hA+SFRzs5Cem6iJWdBd1E4WFo49DCjp1+MENEPYl2xjWxg0hunq7HZtpp7sTesdnztOAxjyNpwGY
upBGWXudgWOpTWNCQzTakDKSjGx4dyw5HwFf2PiDyL/T5tZ59pCcVjpqU/YJi7rxZSJRtpEX1p/o
AEAandKe88h9HzuxILLzvj3yY54Aq8yW6TmYzsijAFqxp1SNcd325Ht5qUBS0m0Aix1GAnXcGprr
7zUqKF91CE6uqJDDoEHns0nJe+5NtxyuQHXBWd4Tw9Pb39eIwygiUHdbAm1Gj7Bj9MmFaWjxmMXW
MgsBuKIyNNx8FZAhHTWRhTk3dld+OlML4ZtrKgpYTAAwzN4I0T38JSXQQYDMteJVp/9XHFZvZdDa
pxyHccKtdGchtYzj7P1PxrXW24W72ZpVZL2upAsDhZph8XL85OoT4lVWpiYySpHvCT4XLBM1aPGb
s+1tqPI3M0KMZScRMZxW95rgMbmJ2bos3v5OZGyUu3OCQqmLL3/WXCxklT241RaYtMhVC0/ONzee
qg2ewzx6tI7aCiv/u4q7Jb4TfwB/t/KZ3akEFU1/nlZx6s1ftebeREEaukakrVIMmOq8l8+OUiUf
EdgoYt07ACucjGpOWVJr/7NPTIuBLg4dj5tb5WlML7G31atX+RDQcG+7YPEBq8i0oozbeLSGo0RQ
lYK2a/hmX0udDMHbaA8S2mrQfVIokxxMm4XVFTadYOjPUWky5oKo53zGHSablYnrJtB4Ky2KRnlg
KqOIVbZzp+ww0uV1KFN7M5ObMBHe8EndBXlfRytvNzByBGmC74eK27WgGN6HrSob6Rn2C3UmQimr
xj+O4MKjMUwuCg70nEcl1wGuhbjNpD9Sl7ZEpIsmIEw+QHvp6H2ndBEWqaASbLLyobelpFw1HzRw
KClqsDTeDog1cPAhoEu8BHRmkddX4zPC7vYtRqDgMXCNIQ20kxt+OEtunr8CfjzBz1VRcWTpC40f
X577mS2FZcC4wuqaNW9FENrkj9ywatD5TGkLg+7oDmiADwyZGeXir+XCay+k2WAi3uwtEyFLyG+K
b1ehqOWcAL9bKtgElclXPkohKvD+QCYB8hoaUJtkV0GG6tyX4SqxAJlAb7lbWTdzuqI0NQrYlxBe
AJjJwDX7uDI7VKxEd2iLq1D9LDgxI2Q3wtDtVHVMcDeaCFpEaeeoE+qry18IAdrfpiwMHMEMT8c6
lSegmyObcZRZlDrWXCLR0B/EOJwfw1Motjz64DFhcHEW2MnREH9haIzdIOGlXFqBIjbjlx+m4TQI
bqMNAGuX4Td7Zqb0BHSG5lAEdAYG+mrR0Jo9L2qntDxWRhuEQt+pcpdG4W5aBzDSoCPjqBNWccLB
7VWcwsF0w0VPGaNYaS19HPvWUf8exNn0zoEYIE4B9eY00wbrfDFqVkw+ZFnGgbuwzBuaw5mfnewT
2WKE1zCLFYj4OOO1KPA0xN54KfxDdPKakWJ+WLFkQwOq2lDYgIFNQZcjGXa1ElnCKYzMYJwqG6sx
xfKWOi77LJsm6kRErboTtNjsi5J0osFo1Uv8eJdR3mMgU6RY6b9ggfpaDITYFjHcKMqMeSRxP3WB
8UIWWR4Dpdsw+QY1wxzgKglKt+kZBmedAhmB7rhHqRni/7qXznxR96jm4KEXJKw+lIbM8hjIjtmh
35qm/pGKdbchGGrq7DdBZnA7WI/JzPTEsLlvER5/vs9qEWqmDRYErUSFcBrA9RE97tAEYKU/qx1U
qBBQSYxJEHF+q1ISBoqIUEak6pWEIEWo+pxD0EIonrH4TqKTOmpxGlWq30r5nwZtdZwlcpdCLkkg
tRYywuf4M+DC4azAMgwvdsu5srm8ah98TX5tq5dp/ACpd1Saq6hjvyJoSTkMYkLu/8uRphCOSeso
Jpax/lais9YJC4yy4hmx6h2rpL/t2VDDK5ynE5aPt76xTdZ/aOlxEKa9SlEPcUsYMlojGbwP5/Wc
bd78CfcUw2wtsEGt9UHSBdlcb/npLQjTjHbeoGdlNhEE82A9wO7mZ+8Ufy0o1m5vbxazj9TT2iBj
Wix1ulnCG3G+b6XmYxZBNLRSQxJdDXDQAvnGqufKfhYKHShV649jTJJOiiwysbOhhh12lyBXocZZ
rPfoWN49QGdQbgRGGg5DRQ+jRE88eb74aZN/kjm3RZGqBEykH9y/KeEEtmxEkgGMXg4bUz2hcXfH
6BSpddy1WGW6AEupbhCT2pXCNtqJkAL4UdY95KA3+R5aNOUw8pHprRzmR0aDyEDGRxS3VrZb+nw8
0KKTlccKJHziuhWtw2fstmDxfS66bgqRvbQARHagnwqmNy8FrQzRquwh5ltrOlmAoSS7McGQslSz
2zco8zs7LtwdIMLY+tjQDgzH293Xwc+B0GuJ4XqK445LP9c8fQe5Fi569cKOJYkKhhkFsPsp294N
+zK1F8QYWrIPoikc0sqpunjAGxbjM0JF8yG4q6FlJuWHuDR/ri9xg0kKnfal1r8R9tNkV5CVCEU3
Ls0jChnT/8uhxkCOitzi7vEfPOj+fap9GIxPPLyl9KZAtemvjgmGU31VTJzjcWwPycYsv3ITgm76
iEGfIIZqXDSQ+vzHEWySt2oXxTnEpSRqEGRyl0zZH2BsWPk58lWQQJbtcgpd4rYHFElMokyvOSeq
trH5Q4vuQOB5/gLPpfcTBpqENhhq5Ecjx5kX9709Bbcchz6IKPQGmPeGgFH3XfFy/CJMOqiFVDb7
zbWlKaXuYxIg8lrILWjh8mDnOgOUzk/o4yQiZSDgl2aUpe/OwOX+34OSeLnOG2vfZBToVCFQfLPU
3lB5e0Fm76WeeWn1zeTOaKFNQWN0uOh9sLyPAaRlyLH2np7lb+OZEhaeAB9WhHVKR3ZTYVZR9L0v
p2q99TQJMZ5bFrsUBpxGm8ASgi0GufusgnqR2nl51sA7ZnMhTPjBdorEVdZgxDnEWv0CK/1gUisG
eEOarRiXc+Nc4/ko5by3xBmgLuLypSxmLFNWbK2UYISZm+NtxAeH1EeZdvWxtgF0Yw9K9jNJMh+i
9D22mwtLNRe2OCRYoYkmOrKzFJZGpACGNp7eAghjEMgopZwnYMLdvIurxhfEGHIq43E0zWoNDln5
gAvHaUtBbHKNdyOYwZ60L2SYXpGxBsXBbHp3PPW6WenFFPWbgav9H3ACTtNjrVykk0WbabYBv8bg
svKrxoj8hdN/JRGNcmr6CKk2fvEX64qTS7sf/OfarzK2v1aAJaGSxkXzMH34B5TxZCeNmJyYRjW5
Q1UAy8xYtE19PuC1N4Ftp6x/JJqh4Y6pTWhmXMfkhX/Blmx1ouv0XRTFek62psYceY+B5B1j/aoM
3Fyd7J7NBIjplBiIQJvJYBxz/PCK4E6bzF7JSU2H3td6HW0ZA34Bxp5kEMLN93uJ6d1OkMEEn87U
cJmmAUzLGqJ4YNhpF69PC+QDKTRCMOVByklFGYzwqC8aaeLHiKiYpfcTKotThp4ijqEo+4cc+hnO
52SVF32zzr3vPlb4J9h1uZmTO3AKpSUrXPcn/KZJTh2IGgbnBWbW6RlVa4uYm9htqdlUN/IYUKUY
N0W7jls3QABk9GYyr3wa1IoEoKpscXhrEQCtymKVrj8KY2shAFZJMq92EeBouR2Ci8JyCv9lP/nO
4fuPgLIjmz1vNJMzKcVEsGEuduezT0BOCrcXXInpDl0XWlYWmXNL2fW3/bpAdVvKJ6izNb6Y+shR
QdZQvGHYFRlM62HCzfO+1oizYaPbweQYXfkEGBO8Klk1aV7GTHJTwhjJNkT+F4wz0/b1oSFzq0a+
9hBZldY5Y2jVGi66EoJxHJyq19/x5DxK0gtrTVc57fv/E+8iAFylcQHXk87nBMKIzSjH6UsztSE/
1ge0XZYBqjwzIdeM2TpGbxs6hgqVpmpj4FySqb0nieyQGsxXxhJQqC6jDlzpVjuAKmvIbIIjs0SH
zHpeilKXLPnz6ZUDgnGvmpUXZbaewzWHLOMWUPTZLW2FmMRSxKffiiqgKDi8CQBt68AcUeRTHudj
Soj/2cL2a54+gCCKn1xUwI1z/ZXtb4Wc052Zjr+wIMXoCzTpCqhb6VEz+zA4rFd9M5qz2jl/ylzR
GDI3lzwVAr1xbMOVzs1m3z3eLydYV582vg58ykyogNnXbeyApJ4PdU2FvFyCou95U0pwfNxpo8f9
sPmBJCOqIWNIr8/TOPgBZF1xBnZWfa6v28KNTR9ZF0CAYZ/DsWA1G0N2X53Xlnk2GiaYq1xzLRB2
0DYUeHXwlpAnlyQ4t+sT96Oxemp8F2ewEVapNwFHXAqLw62qEFe0evC7VCpuEzcNmtN67lWWwnxF
UU1T8Swo9bEBFEvjxmSQxFPv6Fjdf3GFzNRbxZZvtlyJaJ0yox7Ism4jq5ooZdc/8Iy//8C5VEpu
PUypv2r9ZeejAnVy4hDkVbWeHnRcCwTaupU+z5dIOWlGezh5BbVkcbdKH4nGJ8AtbbpCT+DsWjLP
i7krUmIlAQtYU0ibC8oex66X4HOi3L12TU0ZBs0OEK1MDs8KCGfsmOCJeUeTm3P+I39Mt/RLdXod
unoxlTncEKp4JvYnMRR69K2Nwn85bJNX1L12A9A+LCbEp26T0a3Im5IoV0V1DOVWoVUSSqxiJ41Q
KA+pVOqb6HhuLK2vWuHiq6zo52AWbZ/ZIfTNyjz/4kXrhrx01l7DS/AptbFzpvxDf6A81RCHVrgW
4VLaebW5TYjNy/IjoGXc8Sbr3QN1Kndg8K4HUukuIP5H/8a9EFFi8VHVwd+YvUUDvhPm3FnF8twG
jo6G5br4bqyxafco68aqO36zK4cC5dj2LdldF8DEv0R3K100/FPLJ3fXxhD4kIyDDXwfSTMYWkob
y+7d0kGzL27efL6Z0BZ3CCjOIe/4FpC3XbnTeFu8UplblycmMyt9x+qKHxxTCVPAwcuCsKF4iTzT
wDnb1YmtiocEnwBSQyeErupEyEN9S5t+FG6CvuNwXnl+5bp/aaTQuSuHBbBEISN8nxV3K+07KLsJ
b5GSu8UJI/WaIyYQTTuFvkDoksG3QV+3zYku4BrLq8o+C0Oap6QJzmieHpzQeIYnsTmq7uj2fV2F
DobUJ5rZ6s10R2SUuzXGVKJvh8Mh00J5+2Gy4PmCO5OSs3c5ltMjS3WkxUjmHwyUvV/vGhYlZGBM
igBQpRpojpEyekGA9uapfYyNT1Nj55WUWr6qw6uwRB8/fOhFoaJ0ikglXrpUe57rU3KHe9B796J8
O1o7FvXulz0ScIANtvvCixoWfFp3upcJdw1ZlO1f0GE/WUzMcOHCLgAAGmlQChbuBngYGWDACNvL
ppDzXGJd+pZp9djmJXByWFDrZ6LrOdIAe5j42v9dVn+SmkJhUCrY3XdmI0umTJL2jwfGM4lmcj6f
T2Q1K4AGx8oNYOcXVR8OFnB9elNoB6EN7w3EsqpOk/Z+W/2cJKeEAP+O0kEgackwayNd7PJqKoZ1
1NonvPa9hnpsEpeP7JPACXc2tqD1pR3NNDPKYHsCnXVFsgl1pXl/X7kUqttvZsScQ4UZXVy7Od8X
+nBp/JEZ8TpVSy741R5ibzWLEV0cBgbF96sj4gBqv71RrsAxiOplCCo6g7jzjSOIcHc+InHhMJHa
SZlHRfFc/Ftta/ZaHyVnh+RtDA/SEyhPja7nBlRdVLePOuFfOE1MOhzEYsDf3f7JmZlQFLiEegIr
l/9iCUZMUMkpPp2sg7v4k2+xWxVuX/Y7O5ISv0CQbZS7VqrwCm9fvmrdHH3qex8oBpG/OZDRi8vr
OwDYf+NThAn7d+81A1Y2s16p+cNJv6G3BnpZdjZ/JIPsA3YV5ID5DYA+Q+iFNN3gQqSwzyQuZ2uy
EMwhK3s4OJh0Um0Ed7BG9fZ3xxi9INabFJ6z4sMKTZ5Lxqyj6eGd53cP6YZOZeEk9agM8zl4pwRd
tcit4LUqjK3CJQ0Aj7gzQFaBrrZSGRP2bb+AAM1JnGkVIKLVYitBghn1NwwcHqkblwYMdySiWIW0
ZFnkIuNMeLkbqOkwsnPYSiO5SlrcBoqH90k/fscWklFGKHPjD/+v+EJdF/pBy0Eg0ht02+8JxwmM
BbWKET9CPNU6RAl18Z5WK1Yuvl0bkxDSqctsJ73V6wp132AClqwc/Joks17cc/cJ+YwS84LNh7Xx
3mA+ssH+iyAbvvEJJxZeEZQxH6fLrpsZ6Uwifs+0wd+O+ZAWq2BydIfj4dqzSiU2b51MiU1X2c6M
Fylhkc4JPHzSY0MpTykJcOsIx46g1pgdnINg/wIerSrKHaseIw67MWFPhBCWG7lGJl+KeXh9jXVe
hYWkT+wMohDfH8oV6MiRUxA1bE6/nRUEFp5IdpPBLRTusWscpxru3rHa+adtIkGqKBacvpGr+gD5
qurnuws9NzwqN6x5T1T1oYE456/UZhSeRy9tJei0tghkJQELAOaIXsrbQHEIHWqek4XTtdiNnUdq
VqudgjPJUK4+R4iw37Ucm2r72UudJbvVDSRb3bVXu5c6HbS/gwsKShDLaf/ttQdj0RGE36rUw7RQ
0OQxKXfkdTYAfZ6XEl8agx72Vg/Rw/CFsGuXRNaqzJNcZi0H09Ep5jvEhLzB37K6WbkC9LwtNAmR
1cxQ3vit9uhrAluJxqN0VFzFhb766Rpl96h9O2/1VASphNueyhxEuMPiSxNynx4fgKuV1wqX3l9l
kDpOTQ1wCCaE0DzEJq0kSZTQmc8R23LC5AePOD7EaD6vsyDkivxGMfDdFHaBtoLMNSbMTDk6Pmhs
FqRGkbT+5TOH7CQOk3cC8krKuONrzgchp/n08wc/8kM5Ao+ovk5vIYL13hJDHf3I2VuwalOfTfUl
CRIzsgxs5gTjzWwJesYXMmo7K7HKmshSrbVWjiqJoxmJ4R89QJGl/NkCPa0L12ZHWFM2fQ96PPRK
9nyucGlNaC9UYBFGYxFd+JwORDwIPH8LA0RwLkSdKZWIRhE/q9zK0XrrpLXo9aYUXlBHu+9zlp2u
jaSXsF4pAMzKufNpRomtr1YYK4iSGkWYYsxJe5pxCJEc3s9XdNimeH+SfcFCt+ipPxyUxACsds68
ag+ZtfC7vdgNprooRe023RIQ2L+XQ37UIrM4q6o2sEds6oepzJBSwqMn8Xlcr0UPOBrAqRDikyFv
SFh4dtw4W25i0+gvn7cBcWDLumLDC4PQK4L7X4pCe+tZDlTqcAfp+8t+Z9v2ogwBgOJJUwnxjCRN
eJJB+ycbVBIo7iyLo+b+E/6aRbXPOJU69f+2A57ZcikopfQgK+m+t1mGpa/BWpyg1v7md4BvtDuI
burRrC/rAPrVz6s7UXdBWN+dHNsgrcTmOHAGssZ7prVE+W77V6nosmg28p5sUuKF5JebBfk121gG
ykgPmR3+G3k/j/Kfbe9R+POX+uC3EtMky30vvXAZqKCyPvQcyYQP0Q9YpQoq58sIB2sXKDXz78Vi
QQLFpUSxdYEIFzcTaJPPEG6+q90W2nGO8S3ILuMGkYFd4QPmRWAZzCYsgE9Jx2boO1KmN94MJplS
pmMZMJblnhtmMPqUYkHA0JNy+xq3F6QQPDbk9N12MVWY3//hYwIiYcr/FMuMWVQqdzpKmyb0I6Xb
XyI/mO4jGDOQuC+0vzud4g8GHnc12g2c+fZ7ZK+juMyMvyAQr3f92cpAKaTDEKdN4SUSHURM29vT
4Up4/bpHl/XuQkGfrd9d4gRSAK1NaYmbh0KVot6xZ+2k4fZ5Wc9u15DbHm5kyUXwaq0fFRUYB5SM
J025xf+4vwQ7hW6rFvJXr8QGn2MNKEoPuyuvvgx6jonpHTeT6uV7Of6bYdj/9SO2RHjPunEdWwIe
EAr/C/xDxmzxXFEsqKm67dx2CGkUkO4+46910UgRQmS4c9mPUZdfrm1Pgz1TYNTxgkzSragApNKT
ArjEYidsB0TZeKBVobIBM/jiphKcEL+W15dT1D76Mpmzb3wiqniJWUZQozQs+vwYpFGtT/nkCA1f
ySE+kq+8uDF68wIGUqGLZ0tG2KqfFEB09+Yr9gR5m3Fv0JUlXfFAZ4NuBD+LC5N7zOQCk0WhbX00
Un0phX7P6F+i7f3fa7DMkK0NyPIkV2AA7enu0YenrFKUcg/4yP4f3VYxxRMgT7Wep5t4CuXrv6Xh
CHEerJG9fbtZqFaSitCKWf1ib5C+x9FAWcaLkJL6dYhyUG8XlbWJhAYw2bRqeMb6HKAGYZfMyaWT
9F5NAx3OpmObOKq5em8fuq9hhxi9ln2+j8ABr/WTL1abIyjSIjXf/aZgmAJ+nEewhJGICfdNxJ68
CfrTDgqtbMUEaJKKM6KzTXEAw7AlYBczNvGKvtwTCVcr0vf4kFiLj3cVZrH7wYtT/Vmw5Au6yCX3
Nd0I1gbWvG69xEEBZzjnXJA0oVu+mmLpkRZcR+g9oSyGE5lGO4OpOOeln6jOWLPYIMJgw17dIEdl
kwNO/idTpcRiinO7DE0+gNOhw/h6EkFynFdLDFq3eLVp+miYg6P9XCkgV0RVCuVcaYlBaM4vNSof
EXoTtJgGLSWfEcPgS7HzsjoroxKgmQxuqHDkW2BmrA/Tc81IbP1w2vAVmXf6x5GfXSj8YSzM9bSj
aDE5AFe/z3OqKpTOKvvdIQHPuCNPKd43HGCxz+5Qh9h2qa78oQJC05o4bsTHJ7qq0s0FIqEjYH5v
OPKZ9IvFxeQR3aNGSSQzDuSbZ03TtHT067stiWS0obWUGEwZF1Ans128Rcf9/euekDlX8bzGRwrH
FVDFfDsDu071lA/KWBGezbd33/2wjx9R+HugaInlQU5Cq9ATSyd3o/MgEUka7SHkQzWqW6WVn+AH
GlReHW3Cq5u9R2J6csH8G/NzRjSlbDIBHmng44Cl2pRP5X9s8cib8dDCdaEWU3vKYbdPCIvKvPTg
gh2HErLvU4NagL3CLIYHCQlKnGzop+N/v6tH4Q8u3s1VTYv5jvSOcnkH3WFCJXaKqyvs0Geg8jIh
dB9uMzyvECGh47w8w7HLNtd1W7s80TIoAX2iTpVJHBj9hGg8DuTSXEcOXu9b8S5ogh+5t+5jIrcm
0ylh/4ND09qRVd1y6nBxGvS1WexHMkpCLi3gCUdyOrnLGl3dmbIo15q71yD8GpcKRpw8k1rxTXxT
ewjL/+Xhh5eMPmr10ZRjMJspSR+0o8WBPh2KZwVqiPQ2RTsZBgzGqKcPx53Tye4BGDVRRlIhy1ke
FGeaFhuXlLtyONyIFnFkKj+ypBxZYXjhagfkuYOCvNp3QlFGrb3gVU2yMmK56WIxhAumJ142DjUd
RfVT0tk8heMy+abDj2Iap5ac5NpLP7hTj10YZskF44HG5R+ki4f60HKnfX5RxjZlV5WtnHJUWEDO
66izM4F7DH+7lqJtre9YBJeEncpp/OjE+9wwRQRr7hGgRAISNpYOIGi8zgx493b8DEK8G+RF5ZL5
s9UwStJNXKjbY12nco7us+6PnE2fWYRUnRmOOJxj2pVDkoroIgWe77fZN/e7e7JgG4AiU9N44xyb
C33yXIojra47Ap/Dns2CocAw5o/XNyATGyhNu6XQHLYQ2ryjARu5j1Cc2cWqYhDRv3tQE8SZLm+K
hMhLKSdaR3j2upBD8fjOXX3bo10KRg/9ovWa7xA+1aDrdryDdt19LNN7S6VKfu8AYhiudb1q/uOr
QA67KcY9rEhFk4BDGYnfH+54iM+x2D0BdVu3DFxI7Vc1lVYES7HzNSI0o8gw94yJWDMp5m8uvXeM
PPKPhpRWskkNJidyfoQxCbYvXygZSpLfZ9ckcWalmNYY+8fFw2yuFaQAx/FCSs5mIRV7/TLDzfK5
slzozAjCa/F/W6Mh/0S69VwbiMI05Th9G+hoUCDNJHbfQ5MYOfw68rqLjVa3n+lt0cL6GbRRMjKw
FXfJTrQVDjXQXZGu52DrgkoDH2KM3yBPEr8v7V147D1SVT7G+E8DGWqG5HGAU+BWzsdDhZ9hq5y/
c2kEg3rA1n5wJ/iVqwjohHjlcuM1xeqzzCdVXODVO5BLiwj2oYH6UiIW3LC6vDK3NfVAhb27goGE
NRPW78bPK30p8Dz9pb1xwM0uPpCuaikfVGkeKfFp8fHGDBaelFGOfEWI9jBLGnZzAZ3VbZAggDDG
9IMFBhsu1wDDi7Yp56SMp2+bP+FyIuUZ2MnfQfs0asUQBcUtFPU5uO4DqfrrU0DtiedhF87c9/fj
Aq3f8Pm/oztgMvI6m6V+0lG2MnCS+d7R6PPfBs2T6IQ9oLNJnQMvWIaZ2iQHXTbZa9J7NfYvhQLb
TjQoQrXafavLbLUn0ko1cfT3GUnqFakAByo9W/MJkRFozJn8/NYJhCHm6isGJYJ2Q6b4bo3j6mVe
495t8b1MkVo31cYicu4TgVWl2+F71KBVUNytmeaO2030NSo+2Lbinb9Ej4H7/mxs1Vi0G9POrW3Y
h4ma0lm+4Q+sooxZLjB31mla6R21UE9J3flyHjXT19+YRkbZKTI/Hk5g1pPD9MNkssKqId4ltVBx
dIqckIN/mCy3o5IRQC40AOBMXlz57lr5aRo8XKZcdZAgAOEZa8L2J/BLRnX6mI5c6HX4EgMk+Cuu
0m+DLzbebLj+CL6BB7sbqdvO67n/90keJUwDs5T0v5GZl8p2iPT/sRhOUz2FW5FnrKtiFd6f41NS
SLOfZWAQdJRJAkQkjzdMRGQm4zDz7lnxVRaCndRd4LJ6LBDsbjmMl4i/yuPgP+yIAMY8aD7eMkRJ
Jf4IC/fIgm5B7sQIv2Upjrtoozt953IM+oFiZcfSLV87g1woWIYONU3lnxVaEDxzRLGPjBw7J1HF
a5PSxe82NbJ+97KVk7Y4w65VVBrM5bexQM0K/YJishN77kFjIgr1p91n/RiQO3UOSvL2ONGnRPPo
Lv30hZ2gcExRuLJsxI953ddOLRGVXmjLpSgEXMVKFERfwNEblMX3wtGz0jbrFRGKMp8GYoH8Z/Pg
EgSKE5VGLhrlKO4yNC9IunbPko8IqseMvDQI8ZvCLrnlF4Rl8cuVXyCgPRGQayFQhYkpVb/wrOtt
FoRXWYxM6NEvRwAW8HC/jM9KRXh8I7EznxmWqLGrjXY4ypSAl3zOzpAhrWtbHUOZn02WWbG6gUL7
5aCi3Pq5yHRZafFS/bQc6DVSE+1Yit46iWxoxpKm4lFJNI0pWafURGbEblazw0iwH9+upS9vgHbx
Sc7jC2l3df0UHmCMU2PhUSSrAyadzU3cY81PVepLCqbCaSPZb3CvTeeEHYQfPckK7oaP/v5HX35E
0Lkd4r5ZWvVPwsFMORC1e1CpuMQR3BLWtAeTBftYTBwvvcnKtyGSnXyyqaDI4Aato9r/VyvxaPqp
d2Zetq1PtNdGcvem/y8YbasCPbBYgXOE1WeSqzGGZ/L3zPpR7D9qsPNBcKG1pHPbJSNGrcgrKyJa
xSPNBvWlS9EAoKlqZCHa7V5Pwd/PoAIh8Y/2U8lqLJ6fnPN2CG1tPmsD8GMWrYeRJjd73P+rpFub
nHk9U0fNBozC0/puHVxvQrX6srXZ27/AvRTKdE4j6KJvS299eCaORBvV4+hv9qhLq9cSESK9JtiV
cOV5e/slUqnpET9vt+acpuK7YQw+OM/f/gI3cBqLktr3vQkQSTFDBrZpTj7FPVvAmyVgIq4kZ6jS
HJKWM6XB6vV+COOKgtktf+bR4K6upESJmMYFQIaCyTzKDoDOx+k5sB00mALMDc8struJRzVga0ZD
lOh4d7ygpQ78O4kyVtW2wihmdbiri6ck05OJPkIEm1dfRDTn5aSKqjVFaJO0JtFvW0+t4YBQFmI0
MrQEaHyhoq/drqCcZnbScbSGhK8GGMMVNHbJshERZ6DXUEcDRpWkAQVFXYwmRhl/01WgnpCKvpIh
+20HY+SCEVeoeKbf/f/jS/2uqnORZzaygTT4PTWAN6qJaHzSnIshK03i2mKIvztaWej7/xwkzCt0
0bhTFfbCUtDDkrtV83bVpX4z14XCmxi2JsCbhU/SynNOMJsz93fPtrEgLRLcMRMzhbMFbTDfugJO
YPYQAlKpRqdTCyueS+w/UORvbjm9AsAyUaFNlA2J+nAwmzzWlUmSx83ZWmlJG9OL93hXZtXd4c9L
Q5a5Nv0b+z1MCgUQpDe4nTIcWwYl/YXo/V4xInnIbOXeGG/jsBCVJubOIwKzROnNXXQL0SmUsr9w
8cLWqLtLgNo0liyfZbFrbXObv3UeFtasp9HlpwK5n3R1SzaDC2L0cCTudKlXuGZ8Ix1Q9Pa4TRxe
YWfYY14SkcM8pQ2bCrCULZqdI67HyY+6xLAwHiH5lGaOBefajWnmdslIy8UEj+aReOLw9FI4YiZD
RX7yGcYycqy93WAi3SaS7XcVydp8tk8/UzcZDcztMkIaDSvX+ppiwIajM8wbysbPvoZBJKHxoyq3
T8kcw7NabX6O0/l+spTCG0RHozLAEZQyF11Ecvg4Tmi3PXtdHtKeGetpLSDPDyPc8+njhOpcVbak
Gl7/vyj7hBlRacOQKXqMHaO5kW6JNGQWjc7o2RprPG66262jo2hVYeBoufTdSA06iDWb1GLMQOi5
L8q67xE6pB8KsXXljqaroP55nQ5ypK4kujbe6SvVJJTYtkrjfmawrzSNLkutLTmGDJAj75Ui0HDM
4X1V14qv6upa9LltSnSCkJ//61g1xaJW6pRSscVtybUZ2UtmQZ0GDrH/6nk7G9fi6ckw24WplMxM
uWWjc8qAzE3CxpoyEbZkSguLILhmKtF/R7yvWbXgJXr12V609NEU/AtjqvaPo3NlXQR2GCNyph07
Ugq3XZayuqaqB40BA2x4BmcNBrSrYauv1QDealngVA//hYHX+FQ3nwBzBcfl+W8ncL3/NQxCvTgc
L8vBpr4+gg0Kyf5gmyMxV2azf0qJB2nYaxGfTGOjTUajy5J6YGmiZ/EnLjQeK1CNnn/A0dtP9xhm
wJsm/kfa+82vmw4IDdOvhhNB6c7qBZ3WRweVv5TDZUyRNH0JcwUiFvmh47UP1lmgpldzvRDN/KLc
Q11gwA7KJJDx/oyW8YzfMAU5LeVGfHeh0VqdmrQmzxafYCuvapCLC713iDSglh1DdLKS4Rz1d5WB
TWLQlpA9BLXlk8fmmbk67lZewcBl0O4tq5in1PkAl7POEi3IDtT0oO4bprG1KiJv8cqAruecZh+r
eU1azqoA+hUAu//9YWatNLQLGWsaovFNxVwyQyHbS9yHb0lV1dXQuQMkuBbS0/zWasRwUkZRH20u
I+BsmcPkogfUvYwHbjy74ziIRLjiLp4ZDzVyGWmVqXdnnPsFUz3EAWEF4LgptA4cbMl1eiFrvRw/
7H1TTYi+Y+XcVsc1qdk1bFbauwoTGsqYEkCw/psmabvh3QrzgU2IOB1D8yeHOimLD+C60FAOu1QN
teq6MKhlFXlVrsIdyZfduf4fuzwOj2bnDt1/h0j6H9JcOXL59GsbeFtcBVWICb2ZSeHzIYlQQCyu
O2+RxrVRzggNVop2z6d/9QCvOu/posQFXmtCibYYeKyeE//DTYPDrNa3zaIOALI/zkrsmEKNAboW
L3zYXEvEsaAOhAG0rGYIBbXPCzusXR9HnXC/beGRGXNQnLmmJOQuxlAeBSHV679BEiglkA19HUSo
53klFqXPFxphZ8jl18qlx0E35gPCIE3PQGzkovAfP32uww/N8HrFpnWVsnlUKln0+9VcPIr9ftBL
aYHfV9X0dvd7gscJivpdPoxo9WyMcdyJChELSIZnkUHyXyaEnYgXznNqCcba0PZiSdD8sXTdB81K
0E3LInt+kySiT0Cjr8KIH3acTKgq4sme8u/Cuiu8aW6DL7wqtgLPZaf72F91j4TjbS5NkbjbsARI
0YExQKH2ypO/lXbfRWKHm8QVtJrNKImvRpc2LZiv8Hnb0HpkZX7OODbiEYb6+WYIRU62jOy9Kln4
Tt5Jwqls9Rl2PRZHQnoNLj82qlCQGWI7QqUFQw7gciTyOMeIPccuWENnlpXwDSdIgytmWKeLtUOm
2ZtDqKcgH9tcLc7WKMnq+yZ5q7pkkn8A1I9y0BA5HsQf6itHzgDT4GN6UV0vf6Stq38E4xfAvS7u
MvMUGfuCoQE+FMuwisk2o68PpTlsb2qXMbg5MQHkcCbypMmTpBVEMZ9Rv++DzHHM6YfRMP01B+re
nRs4uX+xIPpDW6eSiJyeDzhwQjKq5vVJ0SAKM4RJu2b6Ag1KRvBZ4QxFy4R98Go/vXxL/rlzxF9v
3den3tDrLfj+wLBRiNExYgejDr4w4p61RwfH9DoFhtkWgWVR1E6LS+6B7HMZ+PAzqy9o/UWi2HJE
LmyNffUqEveocNzLGHGeNYL/8tzg4h5jl9wfk4wNJnOz6lBq3/iOj8E2yBN2ZI2lHXfJOFA7oHk1
wOjJ8tYyBq3KbxrvDdAWZLNOfQcYPmLaK47L9lf61r8QP44xPafBuWMFihjzmmWNxeH/O4S04P3d
sbjHJ5nZZkebT06ZZ7sxRYkBjTrfbeuGZ+BPu8kAaNW/HJWC0d/oBpLGAMVRPVgV5roZC8JvYKek
4I4t+3U1hGhjLXfc7v97lefId+FTTNFoTPQAbYTZCHvhs0yfiS3B5k9m3SFOcRugk97P/k+FyfNi
R0pGUfXsTJEQIawvBEd7b204usD6ShsNNEPYcTSBSRdzuPptw7CJLZVZYfGQe55yfsQ5lhh3QYIb
cS4+VrLRoHFdUuz3zAqt0W5ds65hREO8QP45s3/KuoPP6tiPrRnS6QcF+DcFG8G6UtmGVzCMYG6M
LcZF6ufGvZv0CSCdp/C698M3gYvbEe3MTryFwwBn9u7woEbKm/GSbYnGIXSPVYmzcF/hIewmX3wL
VK1ZOxgYS9wc+LW4dSAHBv4g+SFptX21FPw7b1/kM9bUTNpyH6sZkkpU3+5QsON17tQ3eNaEzK5n
3HcoBGL+VPzmye1KSfg9Y1INhTFzifZoubCcufuWUeY1OB5fFCIcHVLujFTM45ocnBWZbehftP8x
dXtzylsuIMvsrdz4ZyYtmC3CJMUfO3dZk+GhkmYR5Gcho6PxZ4xJBIYAkfa+jlak4fRgceJAfR8H
N65MmxW0qPqBMYSrhDX+NEuFZtgmg9YjNo0zQuSLzihLD5vY0Rv0UsORuuK8MNtY9QWBfce0vBfN
+V7hMagJbJo0kQi89AE+aogmjdJJRKhq6aib3ouJXAHrRgSZKOeufSQ90hp7P0DxYEwvkxQpULB7
rN1vNM3i1HuxA5/MNF1LrZ6rKVW1LbYlOQ4d1adlsF5EPN4Pz9Qrv0v923atZvEBneLMEjX/Rv+V
eFPtLYO71UFmVyw31ehotDUgnVzz9gaaBD6+LWhuFkqRljgQY5IWWCHNacW+Mchiq+FyAQsj1J96
bVQOvdEJ65XiQQOkrgyBo/yYX3ve2suL0dcJH3ocTU3qfDoZoT0oNmsv2l1BPY6P7adwjixsv271
XLP1xY3k8xMRhchbzcybXyPHDVddLbKFFp2s+riufxMIJEV4eEAdh0t2JT0SitT/H6YE+z9OAAcN
JSxtozrmCuWal089HMu/3jdrVse68tC1WHveKuq8jnpvziA81JtOGoy5adu1UgjdueSpe5txbOLf
/BAMIY8JqmOlwaNZSIMArHB5oUIMX4bzuuwdksmoxKw65To1Zfx8hXNM5zNCL65BuATOUyrNbMGf
dwiXOn0rPNFcsGAzRPpzJ18klY2FvVe70ldReaUer6xmK1OPENjz1LI7TKPVEI9gpqGN64vbe50H
+xf6nHIg/Xkf16GMbk+awCWTV/ycLB2GV/Yp/9f5N1U+QbjeSPnU//o+0e48qOGXLl4AP3rar8gL
+rTzSTm90zIwsLCUNKm7QuBqXBvl5mZqNjlFwWUMwkSzVufJhfZ3LzWMjlxEm9sLccEmyYF1KKWX
HJj4b0e4jnRheOuh2x/k4CUNY8LtHKUBoVQXEAJsbAL/2zJnphx1SxTRPLEGnIHMmHqnGIVHk1a5
Z/6em9Wn80n1B2GZVqSMXvUG/FmlhoRi9tZbL4S6QTBPkUzDhYQ/WMyzBVMmKRTzMYjUuwp6p3CJ
YdwpB4alW2O2qQhWMXGfI75yqSgLyhRKfW74ZqvYCQwmwH+iNT/VyhufueihULK9NBQYp7PM5WLo
gcKp+I58KlPFsC/qemjNWh9mlIKpZ52nzheO2tXjJiaDklATzOCJs+NGExb80hwB+u4x6ZkClZLL
S1A8KDy2zcmpDz0GJj3ru7ucvyfwc9kddNRGtW2sN7DfkIaDmVymuVMP8atP7SfaTa3ZCCvlCZbz
5Wy++/88vLQ1pIId8SfxUH9rkxMq1hWYfBDctEuONse0oNk9WyD1YB/xV/M4kmmNlT3eQFmlf4Iy
AY5jaEHdkm5SPAQTmUjLIWswiaaFwpYOXLWunh1jZG2OZY+5/tGSw5INiKkMhTwAy1Km17LXKQHR
eIR9/ldvt6lrWRFmPGewYPfw1bSLGFLb+p/p1kJUYP0kAkVHJTZPh7id+AQRaQCPLqlGlF0rK2S6
wEerj4VVl+NNcassWRDSboFWGSAYyMbxdyHokG/o+/CiU68ntpweTCZ3Ds++aNPkjXnT5Mu1KWbH
Ak1deYR8lBx7FrimikMbjn8Z2QVA/v8sRwh2pq4tCTF3SSSzGd26nJ0ybVg+cZEvLUA7PbdldQZf
YkqY0Hwrm9Ypa7YPbnIXJf+QCPqI0kn8XnD08h+mh8THqCuBaxIsFjrW1IqKQThajiUHimvR+CDj
BxJS9XRKa33fyZSd962iqtuoaqBw2GuQ88imQnIOkBk7cgvO6vdBMqoxJqDoTrka1vZzI9vGrTRR
fXEMyVtnDQVsN+jcPNg0FDryn5v98n613lRZ5/8ECYa50hOiNbTm/UY7Smx+kKM1AwZvdAksPNzk
5Ixd1wqndQEnUP775Hod3zq9oez34JWcsVqlShMcScUWVJw106x4cjtaiWIeY8ns4VrL5k+owSlG
oyHihTwQfkEYqvVTCVoYgB89ilcK6gOA7DcwlAEE3RREyXlV9bvla8uaPc4WdAdnReEwo7sVLFK7
YXTfBHXI4fFCDn48ihJEitZi2GGFf3Tv6SAt5EzzKv5/qKEyfp47jv/HojpKux4580BlZLaDTh7R
bOaX004Yn+1kOwfG28KzAGf+2Nx5xsrf8lJyNOaiYygE48eeK5IAVGDcWT1yqhCt/Qi5cCDeHyBg
Z3VjzSjAwBiQIXJVwQ/j/evkd6zrvomGKYXTsOmE1BBPW+oDXUcUg1p1Rq/WahdDb3rh8069swmz
GhKqp3QsVyX80mJ742Ti+Xj0A16adQsSgIu1bofyjEKQCwd4GIyvqofB770jaEGVbCJS61LUPISw
qkSaP3sV8zuEBt1rv7jH4or4prHqbZsKvZ9Cn45WEGPoxbE3YbHQ8ZxtGuPS7pSBakdm+6E1zmb1
n2rRzohC8gHWjmqJGZEQfy2wPgDSPWNEcilPMEmRv1n4Fz9CjtTKEQSQagIMu/Pc4GlOl64YsfO2
nQErmuDQTAWq4/i9aHEuCjT+axM6hGR2LBzmDLXVCdsxmaBJw5YzZpVwSwP/ei0YF9XMEXEP3tIA
nGj0zuP+P5/OIZqwqyRqzA79narAW8SBa7HPOqd9rmX0WRJNo4lsDbX1FlCvOxVMGtYwpwVXp+lA
SaNRxTcbZLJWfT3lIh/w+dOxNgJNcKdnt6hN3C0Mh/Z2psOpiURlEpnp4X3BuLXcwUBK4kQqyQLB
+GirPdSRP5j/3zi7nDLOiPxzfByi6aO7tJNt0MdShjapyxca6PmEu8uN5/M6WfOYu/ugSWA1Jx/b
kr4PB/wna7vix7cpQYt+LuiL7ReZqY229xbmzwkQAsy23MylSDFT/8RUKqeEETudgyLE5yJ6YeUS
jSSNssk6wuGK2UeakxsO3r5kfEBj7FPJwKwaq4Gb/4CFYULwqB9Vwu7WM3ZXlTeMVaMvyPiwIRvY
sNpuCJBSKFPEi9rN+XqM62FYcFY4FLwWoMmIgqY4NOEwHZM+jAUXcTMc0rv2fMzDHYdbyAY41Brm
jtUdMg33D7d1GILAKnvg2iZQapPkdDhyNNEaxuOFNZim05QxvfTfM0YKGqzHGz4QmaX0cLpVa8yy
ClLuooEYBvIVeXrymDC548I7xQExlYv3WzAwq8Qx3aXM8FzQMbFc9qnv0WOuGoUYyfVHRePTa0MY
jXENY7eV7X2rb1txBzDaV9OrasRtMTqw4v3NEtAxxRk1OGgGYWg6gm5twUCOhDbJ68SpsTNY3SE6
kC05qJgwKcGWN5yMalgF5h21UDi/AuY0XmVqB9/409wFZhADBnYN1pTB9xKsCDlxM76mFcp5dwF0
wjzm3+zSQdYUik2S9zaE0ovsvPbc1XP4KJ87FiWcvL0wN0ROtNROIS6xz8b6tPtNaAEla6RH1rGG
N80MbUSB7SB/5iVhqTbtzlxXY1oieJLZ1bXTztz0KuO98ps86B+UbbKWi0D13iIl9qWbL7QdFXSX
edejz7NTkUK/gYkr/ljNMhgDukLAOBYfhyGbmvneS2O8olM+gYh8AeYTjAWrzfFTxqLlCnIEnsQe
THipeFgXAFJHiMApGu9dkvLnlYyQh5k868Lpd7qu6bPoSbU/NWyLWmHC/UcNfnzodm5v6omJnpms
CbDhD0QxOl9+INVyREEjK+BYrXUNVdvZKce9h1GmGjGM8qBg2sI4EOu0lJtoz7wFrnHtguOga/NI
XXQX41SlY1Q8l9nydp7gFVHn39MmTRvg7oqQGCaTiBtqfkxgWFK1ASyrrOC09PvXWdQ2x1loFZCL
ayvSjP8uf+261FXV82lFY6KpjXOGMrd3Gi7zHsDGglZZadViQHKDC6zY+vWnHlNcsCxQGPA5GZij
/lwzErWa21wWGtWFGFxzhLvGFQ22sk6gVU+EyNhtoHY26sJkvINHto0ZKh/0L2pONIVeLKDVfqlW
BA0wrx9lICK3X+zRETBuhEq7BPYcQEsAHsl1YRiS3oAanuyXjQpZgLxPAS5anREGOTkxyNfausOO
V8dz3ikRiExsYvdmyD+cfjFQ051lW3d3dcJbXOLBghkofWCoxbuWsTG8KB2QJLf+6icqrcGL5+pZ
V/QT21f9jk1ZHRz/LZsH1BubM0M7L8SwNj38Ugvrbayr21MFz0FDYfkDL0FX3tKHDrfQTcsLKWyD
mI/tgr1eVE0u7Z01nm3J5hFIucnFLefbWYs+cLQCMdS0Boje5dwt7h7HoTQvTcQPlavqe+CFvHKN
hPPYPITRkGk7J5M8ODkng87soK+xsyklHodHQhX1gp3F2tFE6xzZftmbH4DZCXuiTVitsi1uAWEv
fqIEdMxwqIkWaNjINVOctGPGwRoCWmz8SOmt3WoXX9acsABLr1+xKUJXE+3uX4bMu6OWXD5+f72m
Fy3TKhT0ooJntxsB66k6VH7t/F8G2c/uRNRZuXlOtWdiAZ3ckJ6xvwChJUzOJ1hBrRuaIP1IpJVm
IEgWkVlB+8tP/iRA/X7avGlwuFQm4CCW1e96jwB6HUTCPcc7K0AZvH9khmuR95TtV2FD34/yo3iK
HmsWjb2MKV0XRFO186Q22bNHJCzXxTCTLRVWzctCLADOImTBK7dbIgieikgrizC487fFU4N0tZ2m
bnjdqRs5M2R2ftTFb7mK6cuXOIfeu9tLyD5hn8c0leOgVAlf1j7FMs+KdQMbZjRXZ2Cm4mul6Pl7
ajJCF61kbjl2eAEu26UYxmI9w4Mj/ip1lXCBqv2pBlfEPMYSkV4wlSwiTID5796d7jbkXEBKbKDL
Wh6DPXsIBLMFN+IbSr7BDWNEFTmePS0Yumhuach7gBFpBS7rtBlrosB9SUusfqberLPsCMuIzZsR
m+UDqwvbaoiNlNuiVQ8gKngGsd7mnCHCZdjpwT5ozQUQIGjppqgw1fqHVFgo5dMEAHu+E1Zq2u8u
38A8iks8EV5aExBWD7UdCBj9JoxokCJ/hftIAWn7B7PjzCxLVfkrZWcSIytsBhaelGhgGXw8X6LU
BSk8h9mH42pAX5IYOMtHoqR24btR238HCDHQtpGJ55vBfwb7j9AGoDBrkfvRU9ESl229IuwSLRqi
DgsMO9WYpRryb07OvBmhN0S1SP9DWIlanJzrJCk0+kMVQn8GWSBu+1DrylipfT6k7XzW+d4QWu1L
n/DaR70NyN1Kus5zg26acr15rK7hQyeDD60V6noTV7EnTTIYIHm75BNrqw2os/ErqIcX5zUtNFiB
EYqsGM01SBJ/P+w03K3QWBtlBA82yNwjbuIzuBmHu2dIfzWOC5IoaXphBAdOxsf2argLZp5zMsF9
+QOiHQi9AmZWlLk1Ss6aPOIabXMJKki1uPmkP9+QJ/AWBJvNQSIDl4RmJrMQt29YxICj/0pDhZb3
+MGNdxqQGL8X9xqjLQc47IoXT96TPGSad9GS4v+0vjk+UgjpyriR1PBiyLTfNeWDMwQthceub3bO
bftKLLdptNtJz/1+smq3T0nNX3d04g0RURSEykzyysfxGR5eeiQ/EB+3OsWF3kRtRLantXBCF4Ns
Vr+Ly0UOWwwLxByIEOvCe7CPGmsQZ+mFXknREFMZwKOGsIANG1A5FAsmpy4VWqNH9qtoLYMmJszW
iuz8eyYXO7hAmNBL++pOa7gMl8VmiDDiRP9y3TXErA/SB3tYTouNeS6jTOJCsU52Z2PjwVwgR9z6
lDUGktsUZ0pjVOsd1OzGagYREA4F63Lrvps+s1LXNGzS6fvRavSWfsjV8XPV7FUoHxtYEIjB1c/1
nTIjlgS8/umpCIWfFWa5evPrIbDzJR2wQgcrgp7fTEp0Jl9632zEG57tjGZNwI3Jtdg95/pBnT/8
lduP2UKLqq3eboNcJU8LOaquyCizVE+MXLSBQzRTDyGq/L8eZzhWxYk8sw9BpeZM0dTkIFByTvqv
SszLMdDZX56og8HMoCrI3jLmQhMTxMnMkVZnL0rnz3SzT31MIKUGxGUKqHXxPCF7ooBCJQWoRVzC
eBdAvFfFrZSoc6YrR5qnpGt7oMajM4TYn/dLcg2b5so2431ltZ2QiCzFsd1qqdDesyvFeyIYGNkD
77VFwK/CGSWpPtK+6qxqf/Lp4LYPVu8drqRIJ+COJC4MNx4TEGVLXzGz5EmZr3mvvpZzO6Jx1sxd
o9TmDQqkS2fbAKLzGHpCczG5zT9rsRzqakwB4Ckj6BCIbMsC0GljkyN3B+GGQWEy748pvSe2iTFD
/A09Doogq+6jHl/1FDGJO5G2WyyX3IXShlqyt4KD41O2vAdg4Ua7nO7n1cjyCjAtFLk3+j0vZjaw
kPUhDsFiO6DWCdwapUZVPmzXbxsZOMw/b0+5p02DfthULrZiRB51E+8fE/es5M2934pIxdu5aXS+
jGrOnrMlCA5otph6X11nyN8ngrz5oeTTCJnK7lyLVYqR7i7ezPbx9r0/sTzQxy0aND31DgNbX6ye
lfEqek5bANVayEbcIMsVIgKG8HNcM9rXS3onkjMhPkpwktubPaNi0xEfydkTa3OuYwRyVXsU0OUl
UdLY/I+i4RNkJlRw3lZH6YvkTisGkl3wAJq+lHnT0QpUjEsN7X0zNjfNvI+F3dA5+oCf5+Dnwtdq
QaQ8xcsGuuKhUjTbHiYYR1BzhhEpBqTBMVfLZintuw/YOx/0LADnwu0yPtsKohGUuTfHQRYN+oQH
3YnduSDCKl4uuaWHFi9acZQ0+I2hZhuTUAIvnLel6nWoNB2TNM+9eM57Na4o6h1wmFr5LWOAYng3
9NAHpvJlYo68vLbWuKz6piDrdq54GGnAlrh8chzWVjl8pIy/N8NcIWZVUZBGTVof0DiCC3k6TxRx
P8gBdVt0ssT54+o+dDKp38RrlHr6fPcShP1fBhjaFb5OyeIBNzs31ynNOm61uV9iPBZAXjjm1/+v
3FV4yKOAyqZUwatiBM1gFKvhxpaXF8LYBu2i0pgUwdW+dLwfQalkXUJM/iBDJIfAGIMyhpsdBISM
H2Y4V3VIc2gN5I89uW6jY5fIjMALnDwzMTy8OCEZIg/L93fPBG10vzwSFEYVk9TkZGQiRCfyjUH/
Q0et24aLmZHlGQV4Jr50x38LApWYS302mIjSlr64q1qFK6rYWQewQUe48R80DpIEAbV0d52cf1Sv
r98JJlDds0WStSc2G0USu5oQCatSzA6NTyMx6jjLg3R2kTPR+GIb7O2C23rqdGZ+jDWFH8QIG+XY
XYu50AM88+/pW45PqN2Th4q2R4hflwvcDu4NIua+doDEY0bzwc+79OAhkos77IPtfgxTiQAKfaw1
g7Mfx97zeUtef/Aabj9pSJmiiov0vwXVACH16b+DqWUOlde4I2ocNAMta9XVQsU3vE+SWu/EuaTK
mry6uUjfl2jGKJazeeOFZUmyh8vcHcp0/9HgLaes3I0Esizu12NFqrkovqpHj4zUkvL+UvSxne34
zWDHGlELxCflsM3fBj1p5MiGYmjY+XWUo3tQagziYS38SbhazzIRP8jWZ1Y1LdzAAidbFIpRw8g/
E/IRP+GcrsuJS4jkKgFcRTo/cvuzPcHaXieg4rNRL8QZPAJf8hirAo2/1JD+5ZgmWfXM7hdllrxZ
9rQYBC2nNZ1mNklVclk9t3ryga20MVvJCJ5k7cSHBfo+eNmrwz+Fjfp0D5P34ZN4mSacg4shhvKa
YWfAzAnMTGYkhMz9F9DeixY0d37P0uSw+j++VjFZkR5hBXSDES4ZtAg8sfcGAnlq0fUqVyOO+CHM
dpzYJDJvad2hKhV++CXgPHqKUl6mRdpv9fHERLBLCaz+DqnkQuMrKZoNo7fb5NtJiSTyf3nV9bb/
2ATNAfBnh6T/4pI4J2ri+57KLRDRq8yRQx+ZaaVBZs6QWhTmASX2/HjKV1k4GpqnFsImceyiXLIH
bfLXE07NupZJw9IX/e9sixEr/BLMI8f+wRTiQD9ls7HAReaJQeYVz9dNHfXU0P0mwI+S/OqBmqPu
EEe4p4vFoHGcXVcVA+I2Suoh9QTOovDJ32saMizTash0EhQ8pYVQiVIekAVafb3jIuBfD/ARfELC
+4A/DtHd60FNQIbFKWQyHZ6+qlGf0ug2wKcgz0wdykyZHeRKluvz7pyfE1tvqgMgFzXriPYC4WNG
8I9k7yvKRGj9U11LRIuNQNa6HCorKm9zzUOMV3Wpwc6apcOaMYANpib3y+wPl2kmJ3B14Ws9wTGN
up+l41JHPiluJ3QgdTgr4nIp/7MFWZsTmBRhqOxfgrlfX30UrQZ1aKoTGPeVMZd7TbKn8BsJBSDa
RPTegLt/abWVcgzo33oAYqvfFseGzqrgTOZBixBv0S2LNSvBtzu1gY584BZfIW484Kn1Q8SC3YJi
/y+YBFNY6aB2f1R0yfYRa5GbVbuPwm6pSgzeuOOdbPNk+FTugooNldwUfLNUWdjuyrykgLhdyLXP
pYzkK/Rpv5aI8QT7LlPi3Tul1Epv16JzFik26NhyC52VBcm3HbJVX6PZ+dCtGwIjLhdW2mQ/eXiG
iLt1t761KjNMRsEkdd5mIvqXW8DHh4Yucl/TVNrdjF+6RFgXd5An4H/qBc9jVHyboHjnFR7j7pgx
0exOYd8qOtAYHV6td8udO15dGMIGKX2LlyqQQi0T5VXgg/BQhZnLhXvgoeeK3892BuJZetG7xWfW
GKGGVAsvYpVa+Q1XhGha5DU+IAicaN7SNn4Z4JnxHv8bh8r9G8Voee22b5oAp3vYTNg/KBxCRcBZ
rPEeCYBjR+MKhWuz2zecYp5AbncsE9wBQY3fPS0N9mqidZDtGxZQiY0AZvkr12i7cKj6iqcqe0pv
CgjBWMYu42vMjHj6hFm0LYBmsHQvV+4eW8WnKoIulzJfO1RkpxnplEskdZYrLSh0WZAwKv8LjU8W
ctQl8VyFz/jVMjXIka49qSirXBb2u7au9InShPIGI1ZfKFIjEYdJtk+LxflQDCFg7QmUBt7E9uRu
B/KqiYRwgkcWr1ugiPe2GgiZnj2lUdWysv9gzHVqICO4ZHjDZLAQs1DFXCgWDdTShPWxcoDQDrHW
0qNQ0frNxA7h8DHeCGG9vdZFvLspPaxryrwPbjxgVZZNecO7F8Y0+nkyXMMg73TSJzIb2NFyIR7D
0U2l1XsUhswnEMl7cB9eUv0nKE8whHUfg+ky1pwEfGIQpF2gFcV43wsXfERjesAUYaQJGGmfQCZG
j9o9gMXpw2CcqZWbQmqHusxWIGstsF2ecIsYQdFRozQtC8foDFf0Ul1LJLUKTsfNWeG1qOl8kmZX
d8QrJ/7EmddRhhKxkC6+1o6sGZrBmQqajKWE22y9HNLEXtwMMwvuE+3ywD5qiIYHdZE8W6k4377z
onOrzCkobY2bIa4hkLHbISSiwxLmmEE5ue/T/LhRsS6kdABy9L86J7T4d26K0kVl8hn0NxSJ/NVb
TSNI60JQZmINhvNM2L3FoK1kBbSDu6IqdRVZ577P5VpEd2Dn0tSdUPyqTncbHmV568BXWzlsdogv
yNnyQ4PLFyjkpNiKmNpmFx2vbQL0GgRUR5qsxyOkumKgTFQrGN/AQQPecAmvyyX1xHedT+fYJCRG
VoViJeSPtBv9V35KfiLO0zNB9v8EGzTeqDcg9Dn71AgyTbwo0FEEAiLfs12IdGXOYsnLiHWkR+vr
m5oYTYTGf+F/IRUcqF01dYnoWRVWmA3TkOy2ANSAC5FamF8rI4dq+QDAcJe6NbTpmkpEgtIjtx79
tB2C3/6YhC1dw+6kS6HbNcAxywia38+C2pJNmPH5zmUh/VxtunaALGwpCMKZEsbafM62zZo1HXSF
kYlrMRL6HUxY1UyE74pb2brzC83OZCJqUfPmdiU0zd2z0D0Wx2zViQclQur7QMiUWTT/d/o6iN3M
l8PzaB3Mrd+GWY0cLhcyqAeUs8kKI3y8215vwUoBAQC3bb8nAuj5584wK4B6Za0NUa+yv9dGx+DX
bs4VU9rqS9zntSjndXHcn7dxlTQ5/FHxxri7vAcY86i0Ibw0LIl5iaPWb+Cy5/ieftwUqxWW5O8O
58W1FVzdnqReifncGI1pjOqpnWzVM8lea+97MC6PqsusuFkcz0TAd+qow2MFpqmqxwo+IHzCfyTk
igE7IKZzwY2dNIb6tICHeSVx+D4gO8oiU9Fsq7OWgPaJ0lUxGQK4CWyW61qmphwPEP+Tx+RiJgBr
pjuLVMUfMMNGBlQyuDC6yRVdb4Ua5loXG9/2k7dfPQPSinhD6rjQgxbhppFu7wVPNrMgXD3tfpih
Jbqa/Hk9RMcB84dwdan78nRNz881tNs56Pn9bNOtQjiEsmSHOfrtSplLoAh3JEZFOjLjMB/BmEll
YuBuarFXF+ECNZlE22k/weLf58D3cDRimo/hicS6ne7646hrAdTpubTUNi9DYBnh6386EKkOFCiV
SljGVZc4MNIhjDk2lEPoZP8Y3yrjneiPy5b7rXoOw/aJE1zaeSkvtWOvFQ0hKpbWHDPWnkM1EzRu
rQPJNqzGjFhg5Yhm6g6pG5qTTufjDCPBZYy4R/nAgQwqXad3qYzX1oqQrJxaKjjAf0mlJ3SSsAUE
zC3oBjrYHO7lgoAxRLfaI+BGC3FF9XA8u0U3RYzEm3hx4I/jWRiVukIcrTigBztWHVz016k7SwG7
EzhlCtr6Qpulcc57icix0buGmT/GWnqDNwgfQS3jBbHHg96DvE6m83UKqUrlsY8bNKMWE6giZ/t8
BXrTjtdJVd7Lw+VNS3v8Cw4/wl/ODjqp5n06pKYi6SfKj4bDEgPG1A87KUdnQMe8fU5A7nwQdU5v
f0+SKwZDqqII2pVXaK7Lh1bF5nfVRSaWXWa8GJoE2RNpT3bKKRLHkwqMbw527VmjRwFoHT79kblc
GHDo/E8D7kwIL+GXSuoA9TtMiQowSlULi5+NoiNy+hbk14LkgQBbK7FIGg7KCntYnB+/IdN9ePJm
+FwzgWHKRBWgwllSWki6oEO6SuWu7YQRt0AqrY9auCJdaG2t4aVjBt0lBnNJEPiaO1bCAZoqhV4H
UJ1KBVm1P1LDHF6wm5XrbICBoiUshke4mui6dSicxt0wwn2J4X5tUD7K4LZ0CnVrCiQ9rnf25f06
zveoG0IliAJSNu2GJiJlB0iJHt3HaTaI9A3Ja5STgPAyMXch3xmnJYbHPvG154iGHTGdcabyIQxE
oafmqnH0PdDCfFy2ivHd+NMobOtbyLrapX/bQuMUghxchEcuCoGWtUOtWAbgxn1rkzHsjwbilrIN
t1dcVnxQHuFeGDdZWwFPV0JZ9S6maL5KcQf7j1aPIJYWtWFzfMYo2dZfrun7hZlwoGWShWi7/2eT
MWED7yR8t7UVxXvnXHZOTVqTaU5p+HmrPmwmJIz2O6Cf4bX0M4M9Vok8D7Gdy5qICVO5QtKptKz8
QhTb9mKV9sI6rmHPBRjW0/UZYYkGao8j4akaGLKkwkqubpx3R+61C4VfloMb/FxErGN08KymgcRF
r91TmC/zJZOlOkANsfkRmjpP8u/zz5YNbZl4kj1ms02N5Q+hi6m6rS8S03NHAvSoSTQCGcYLs8jJ
1JZERmIhpTSfW692Hr/Ku7K65SbkA2KMR+Yq9+hNjXVy0L34kjwxoIQ88w6r8I5/HLCB0zd8cQp5
9K1RadfAA94i2O/cna/e46gpdwen7mKvHbgveZY7J/VkCBhShvrpAxpkqurWCDd2XKkjRNzf34it
ChSFxjhM+PSW0URQSHvUslpaqb89aOVj9MFoYvOtII6w65I6SSUEr+BXfflpaY5Y5uMwzRKgxsDj
ggN27vD2EAd8mCJuYq8euu5eqwPINq6um0rDrXWUIpXyqe6frmrJpXWmpZfif+M5oR6MJBUtN8U7
oSaEmB5L4k0yXBjbJw1tq74SwDAEhRGdvVJP9xJTYUhoz95YOOjkcPvDAo1sMQ/mUWUhrC1M/Ckd
DgWw0lfQi4S9Qu4Tf6rrR8F0TDvGJ4F/aTlhgz4Hdj/nfyHP2tFco31/i1KLcipov4VOVByQekuk
fJDW5eWnpExCKrZjyFZlu0xnD57LNmNYCOkdusmdHwUY3UtaX+uJff+Yz/gWc5cV1kw9IGHuVUa/
Bc4io8/Kl9WppECNxH55XQKgS0W/PCcOTQkg2a92UO5M8YLvTG85a6E7cstYMLVvADExDr3Xnqn3
Xi9kLktFlBJcU+4JxC9epn1NJCOQg4SXK7P1baJOiZXVnPMFe0rePVyLoc6bVANJOg3M/0KubEv6
1ZE6uKaX9zXgKKt1Rta4BxTahypW9SCN/Ufqm/R5/9hdweiD0lYt50O62AIkP705KJIY7QxrFUVX
w2bB8VX+DNo+NTrN7eHscYPIYXd2zx8HgfO4Td4Wxd2I8szpkM7q+gVwfrBw1P3SCfR//5K5QWFr
guqz3CHQ8Tmdh8dikDPI9PptuYZEupt5FD/xjWSTr0B7Tl5Ftmx0lpyYJEClvh/Ye7NVFR2s+9pd
oRu5cNE6VfK62zLLqUXmhb5ISlc0+sryw4j5jAGOJOnLjnRmMUx6ARTndzSokV5lTQM/qX2VvWLh
PUHscR8S2s4EZGeUSlzpPUWSiEV1+NIPk2GajuHU722f5nFm8aWK36cf7Paq3JfgTzTobFPB08J3
/1tV1rnfz1rLrENk4Xx1mx4tVY83cL8EaQWZJDYikck/h2ieAIv5hCatpL4if1D3VldjsK/mPf6/
1k1ogar0nXJi4/WPcUf96J1MJkw4iBwefco2Oo0qnM24wbmUS/BRyUN+vaVKWSmc5MZlBzEBNm99
HfJQxmIwGYYk4FJlNNOnauEniuFahjpFCE6k4ANiz4yPY205ubR83ZmtiNAc17AwuQxwIdFemLDG
NIhfji/ne9EVQhIoHaIDLlufm+fRgVwrGjJUTULmOWxzE3wOJxDkYxO/JnqFj5SS7Dg6XLHKsfgF
kgD2iZReW5Fej501Yy9AELS60yvmze0DzRzmvwUahNogoJL9LeubBhwReQDX+G6cZmiDJzM3a0CU
SxCe1AxxKKoN4OFisVpxCuTs/bqo4nL1Y0O4YhguOGT9s610poH0TRDRMcpuNeLnw12unXrdwFHI
ZRzYEUjSc7XB6Pl14NQkc8xmUM4mPkz0nUQI3y49KaD79ep1jqyfS/psRp4c2XnY9ZS5Ld6VRyXx
JkMW32rLMtKWhTvIPP9XWkcK64MOJ+jLr0Py2+SJLf6DWnOCWVKaGX0Jaftx7glfx403GmzXQ8hz
NXiMRzEu3d+5C4F0Ap7lU62vch3ahaiJojBM+98+EsVrF3V+4cDAMFfqjuqYfqdwfz/yDF1Qi/Mr
A14qExJv7sOkR48dxVBl6gBvJE/AgdmYCrXDE8MZatAAMTB2Rj0IFKhHy/ve7d8OOW7+kdXHnxce
D+d63WA3Y/AGQxq3fBXcGJqwCcP94s8CyZI1b/R3di2mFH1dbjfF/6SwHeflatwu8c/Z7fdDzaSr
tSx/LR2Lw6gO85ssdEZow3bVhUA3D1CXVWmCMHRa2PwuxltseQDoIBNlQQN7QdO93hheS+9Brrv+
IhI3Yb1JBvuoO+6/L3/tNR9lsAo5C4rXTB1nX5idyJCWYT4q9s9LjWOuQr0RwaPxXGrzYyQ9gCBe
QVdmFmtl3ntNsWlLwhnwxty7EidSg/ovibAqabBnRzelJ93XoABSSY7shhV2T0k0QbUGfK9jQ9oc
HXRixVuhY4ENzGz62g2NUYiojHFWAqbQuNYRD/0r74/pVA90xG+7/eTxDN3lpSjXGVGpJy+5ZCOa
wpIJl8InbtY1810ebCgjslqTgPjmRu0JGebKwopXTp8qqXUew9rlq/EsTZNuYPr75QcJNkduOyoW
coqMnet+i5vcuP6ZVYCJl60usHNZXTZwls5e7yHUjOiouN8GavmSO1jRvqyt6YUdviFyWCD4Xe/B
aLmaWBQx0LGU4wc5y6GFHpfyZvc4h54cz1+R4xtd9GzNuVgHmDerBeOX11GpeBD1ZkxexHDBc0Pp
HiHU9hrMH2pr4bCfJonstySu0Zu4Vr90JLuEQJoklveyuhQRAr2NY79m4jbYq0DhNe2qK42XzYsH
i0ZCMYoMyVWRaRFJu8pYGKF6SKE/M1SXWEYHEPIaF3tkkTJKVBIn6LgTiVY5djpsYaKEOE9j3N61
tPNIpc4vhrMOJgQaSh3hrlv2Khhf5yjWXdW8Ys+YONawkOAxhwGkrJrfS/GU0rVb3w/tUrywkA56
jiLyAju4xngKrlskMlxpzylYLDEe4up3/7c0/9j97ZLnodX5uuh4S+QHGPYuz4V4JUq2y7kU1rDt
u4/D0s3P/BQPPRWtBl2q9A0nr+RANpfQ0HeT83V0G0NMUEorI0F6CkKD1yEYDkltqPemx0uz0bPf
P6+BjsLFfzeMabqFZ5MxBQGBeZBnlRyyeOFmGwpznNfaj/JunaQERBBmym3jgs26XFcgMc5pV465
W4bWSXnJ6dKeZLB9jDn2cZkM66QM47VrhI53BQoPtbHZfOTmXDsEGanlgsZ7GSoTP0oNCsXf0PAu
oCZxKTcx+Cu3xLs9ZpfiVIPJ/YqhsN/KM64WLq516TKB7BTMqF1nKcx3i3EvD+i6/6aNlv/sj9Lg
6+KMcTNqTdOJahtCxZj9IW+iJyFWEe3EfNj8ZMmmsrbXk7i9fKQUGvY019tCEhZjioiytEC7Jn6j
jU71HKyN6XahHdgaeOIubIh372+lKZL29svQwAlqOtjamY2E/FSHks209m+vmpmSO19ahcXufCnN
bdAfAIpFGF6r5WerdVhcdbMD+XxxyajkCy1buTNYXOszewpwrK5i41hITKUjdvmUOxCb9nute7OC
OnmXqr76b52ctOmmpyKh/7Lrr99s4d6XA4X8IL84wk9a/f4u7jm7EudBRaCXgus8JaPifEdPHRJh
oJtbgFiLToRNJn4N3xMa3ASAdojZk90NhBkIEmpY3LvfZXwtFyTXmG6Xbd6JfkN8XFitaiGd+1PM
qZTZXL+zlN0c2AnY1zPTT+haROXzAn3NBY2nVAq7dwlIycoBOvzDJL3Vah1QP4FmvBJ2TGdpPNZw
Bbgi5AG8x0VG/Ke+YqXEutzCdlXTVhTpDbYGdg9M8Iy5519kSf1ppNPjUcZVhE0eTfZHvbHau/kW
urhEMfVOr4v/ggwhoneJ1dfCVucd3gt+ixISAtoKtselp66n+7VZIW3DsDHXOFJj1+pMmjjcd0F5
UaiaWCv7wPjoQSAlL4/3UqV/75fUhhpjxa/zx1aqJ3C1E7dCMz3SulhvqYAVB4r2BjJvQprzhFRr
tNxv/PNG9qbhUz77Bfb0svXfyNNtQpiBLGaWb9K8mZLa16Nd6NcGHfdj9kOto1qXvizIeYZlRr0o
Xv45BDDebEit5dfr1kGWlavh4cGqYm5MUSvUYqLRv0VY5EiWbTx/7KzTQcKuP9QWOv/MxYp3AzYa
oF5dsuimve+zW0FzlojYAov8NudXCPAcC8dPvQ+dFBUQtHbzRtQbZ94j4/GEGyQbvahK2PtjpkoI
l00xtWQ8xfxnQ5zKC+Mpx60vk8mpmxSKIIW0DksqtBBxUXRzjOrG3NZXpFdYIkcwJVBmRkwwEURZ
5IsTyBXUU8ImSLBOhv2OtVPrrmfu/RjFCvEKzOcjcitCe4Hrj7k6RbEd73F8xw2gbgzEv97D5yiU
p1wmtRX9k4HOiOJg9vUq76DBkq6fAgzedgHQScrTM/smCbK0tTo85730hyZlyK8hyo8vplnu9/GB
UTrZiBFN9uZWL0L5PQiW5bSiYHP9JgUzgGwrrZ/z+FupgZRLYiZF5OkLaVd2ayzKEdE6rd73X7QX
qvwXr1yVsVL6fYUZXI2TnkZOl/DmvkXTCOekMr7QyVWHdMnSAd/69+9ENtfOkwVqaB6EFOjJCWMr
bb1eTj/YLJa/agF+G3cRMu5QksLdGSUnr8ukShnmmcxLWMSEsRjPqVBhg7cAVNdkuKp7nYj22cZ/
xHM3uOL3JQYsY2zQNa92xL4IOf7QUMyPnuk7baP/FsUqUrk6EYJ5sOI4f3fEIqSX4rMHVKwbNj3m
G++TLJ2E7NFz3dr6hxrOhn3EOFM/lctdN2mAr15Ql/EyAyBH3CoB1MYWh5OdQXiFxLqXNKOn3fgR
Nv375DC3YQp73sSzFq8zPAMvMKzTqt/wZ0uly0PU4qiwg0q5SpLT9jzgjqo/Q1bzxe9uaQ39SHk6
KYe3mVBhFdqpzOjXSS27ABisRUPDhZe+M453Bmv9RKXaGCNgSAIe9Bvey5bMeH+VPBnex3VgavSf
NKeDjjyVWtU5+3WjxkMT8JWOhmnSYnP6sZztTxA8MWUjMEnl8HuFlddmUKq2i3ipCjL75VVmzAiN
ICsKnaGlgtMeDSZavYJ46zjuhsOFcQOYtUS0RFyyw9Shv1xUdbcbn1W6xdaHANwUM7J20POzu+1i
BQ9Ikho35RjQYaPW5bWSy8BPjbFsE/WGtQGTYsw3ypwUolSndmhrsvTi+hvU4qV7In2Q/5/jcEvt
37T2JOoNgss5qxoUWZxRzwU5o+4TVMrVe4YqVw3hch68sriFFzZJUn6CVXn/rT5fxWnU8NC1GLK0
6wObUNMy014qmzZ9p8gjnPWgNuo+RQ6W70uFNuHyckFuc8PS9VjiW0smmFUgNxjCj8rphJRmUqfG
xqD7cpbrd9qws/bYW/X6YNNifpy4RnntxLhP4fTFGuHqjQm6MVwH3eej348oRRGdek/FuQFBetYd
GcQGQjJCovI6SRE7prnqtrs3sy2KF7MoLwrQuhxPd6LTekYou5aSNE0Xqu0JjCwE5z2BuKQiK14g
4B9vx8iKMQ0iVypzsDBn+p9bTuTwP2Wc2l+S2kU9x2fttqD/xP7LYEKJ8o8/w2uDfDop4N/bZbqn
lZ+nzVgwI5IuwIAs/VfMr8g+xwgX7+2M7WTLV6hqB/pf7PLeMfZ997CmkAjRDKfT/zmfDCR3V42k
Py79N3FGpPMIgY4q9nA8hGy4junjebtd+1sDTZp1yCt9Nc1aW0LiOvFDTIhUSj9h25U8/FP66V6z
grlAFuKCmM95qhJmfCYHEbQeblGxJfB5Zr+YJxzBvS4RQrD45h7Y2BKlVUbGHhJFnUyOPW0QE8fX
ZM9z0SlDjgmzv+2VA2PkmJK4QMcUuwA4lCHRTJO3FWM9swAgN6gfPUVfejRqg+M/DPfryxgeZDwJ
bHCrc2+62iNIr28Yfu1EuVpoU4TyODw0ehD5hynrraGQ9UcP24NDEiinNPrrnQWk85UypaBz6KMU
g/M00IXq1wLCUuoNGklWcWxd1/HJoHYf77POtZ4Fw/3mLGXvsUrX9gZwI6N3pK2GwJT8ThA9/MQf
lGVsbOeJq2ndPMcl5iH9MfGnBv2GQveNcQJ8MxLv+QMmWwQV/2pAYaHwAWp+P+YW22yUlTvycmR0
a/1IXu4y7z5B/UdFEg8aQMW85FI97/TNgppFigP9jdUIf/cDO6Qy69H8JmUkYvEDl6CvSKZPdPxy
GFwy+yG4XY/POVfwrvsvwMpX7a95ifOQ+j0yoz8cAeI2gRSHTZpj3Npd+ThT2i+DNGhZUcEJkBGM
Krdv98UW1AY9B0WPtu/kCegapfEzd3SiRR0zOdOZ4wLqZIKUmuzqhLQBQKKtsRt7V4E2+ZXSg0rQ
IaS37XmLS3nFsY+yKbxiN1Kwkz7GSHD4ouTr/jfvUpWntkzAk+yhZEi3IIdxyOKki0b/AmfSEqOb
sxFyIKjNm+XWaSXDjS8dzoBegVBSR40tShip03TUZHD/BOLYa4jwKqsIdWqpe8X6b/OFXqyvY6Y9
dpDkLLBX9vIFGcKxbLWW9gUkzdgKSZAWZO+YFrXchTvPvrrczrH2sFhj+jPtXQmBAKh1448G5AWv
DnNiXN2Kdg9GC5TIFxdyQcDSUnF4jGq4IdmWRMmkdHZ5jmETd/OK1N5PhhBgOTjbiNXLU4uXnCbL
yr8lq+NWHOu/FFQEYYzQKFCnWmvsn/TiFnFztKbsb9ZophDkOuE14Yz7CKge9I8EOFpyUIm+GxvZ
9DVaPpmKoINiy13MsAXIYpaL17tgaX/oahNMZ4Uqy3eWByLq2Wv0Y90rQKzsd8RQOYEpW/jDwGsS
5GIOwv0j7OeZ7snHG8by78u9wF5mcyVTOutkTgo07eTpZR+DYpHeTbPbjxfIO2zb79Cmu61hZR83
fWVr8OpdZhkGvvBeE0zmpVpp+KcmY84tqwroeXuDIJffZAVvdqsAM/6BDdhR08i4CclzMXuhVeyQ
mIiemeom6/BGKMHBjeix5wPRRijeJY4L2kwE7gN7UfDnOF2OIVhvEZQeXsx/5ikhH4reiucGmH6A
ytSW6XUpAZGR/btx9QfEUHbKVfMf73xfAfelDrj2SK5KXIFYf/dNXhc/56tqcz71nQTBrTDqqRX8
zMWQMZquviodzs2YWtXFykeBe3wTt/nUeVQPUcS3bBbYtvf3We6/u3dme7MytZUWZyDn6YTrE50R
ydVjs3uV55vyVXONeK1sC1Fc8BtLGt2P+bY4Zu/0op9kAwo4fWCusDxtrk6M0lDgGh6prKeFMBB9
EydJJCLUi/SZaWGM+1SG+VUOxNAwTCjqisIbR5JGqBhde8FfppFLkZG7Rq7p/gerqEYrV61KwowX
P8KsalDW+wkTyq4WGiVgAeVgD1HNCtzt0rOJD229JE8/o76HD+NaTZlWL6XBN/w3+p9vqv6yu9to
gjJA4+xCInKLSVUSzenbIJfVvtRFTCY+HvkdTK0iS9TzXxetDag+ITtPPFgxKz0ybSPDGRKv+Wju
0MFIumuhpDSPYDIFtgZq813RrQUzV8dXRtE+qAMA2fWr3xZciftPOvbfVsBlkQ3YqytaClqvKOmd
yjPLwuhI5ZimBxcvyt2ZTnOa8B8JlBCZWFHZuYxOeG0dBezKOkzVXhstTL3i4XRNG5om94iOcenj
7/4DEeGCO765ymd398kMBdS/pKOPdNS0u28P1C2rnJog40sA0/46bgKziwLeu1+ZplzcKe58EwZQ
My/2UGk3E3EsiCn/4Reu9qTSjmA6TLybwVEAKERZKOB5eb+lYp/rjnBP+6kV3++Y14qQS4pnCCE/
N9sfbT+jAo0vvmm9AufY5h1vdMRHl98nzvsS8bXouaP39fmd3ecc5ZI6j1B6qJ+heU5iTA/azJDT
ZL1BdTgMpTCOLAZzsiwkgaJzcTq4O0u+wYuhHXqi4dcWT24Gvf9K4ac2/uM/JYV3SHE3kxT5pO8K
obX9Rlm6eZJAmIA/Crj2WIP7xCcky07ByQdFg6+y41dxheAT9UrwFiTeb5uGHBo1la6kvHlj7Dh2
RR1XJE+AZLs923nYWQHxo52ZZt6tfE7D49Rm+PAs5nRTacn7DBEaTW7YZTMdkcXEnr+5XmXVwEow
IT38EcuFNpc+1bIRktCE1uwtaH2y3Xwe1WHWcBhKz9Bf6q7LpS5PqeeNJgov8EJMI5DFYZUdyIYh
3jAJ3pNTIctxPObLL5ymJewtU+bAmyo+PG/pirat26c6R59ywzYJoYw7o9xX6nZw0BUHEQ2Or8k1
UdcfyDSkRzpJkTMWBfqowPl7owxIIU/MnJCofwj+CPfhkMxvN75fMOFg6j8AY0Ffi/FocLio6ANQ
AakWvCSiV+TQWGoYObHJBqHrid+T6I6Vc0zg+gCgaKq/H7OKBPpPU3yUQ5M4uGnfGxCrWW3/JYlj
gnCeNg6Y9e47xUP9Inve2V0pcTCCZxp0KMgSqA6Vd94+KZ+yMZU1AdzGjhurQF2N/PvuspFGYnnv
0tnEqUpogrm4ogRAZ/G+cbK8hR4nugtQXuUV2CEJFcSX8wWVth/dQU4e4kowZgeHQG3BR5xbfmSZ
nKz6lMg5qtpM0yD8z2tsKFB9Ywc03qEwpmdGq2FhQYJbTTWTgh7wvnWiCIyU3ZzINeGsHsA9IIoO
C4iuK7z9ZD4g0jFmS2SlhS43IQcWd1kYhXo6kjOpM6QzPJxuHg7r4ZpUkCQcCglAoWbjUu2uPbVe
PFeNIebhS6uz3ElYE8WSmI8XxrbLx0e7wYaxYxNI7i6iEUSDS7GEEOO5Lb+ELjNgIm6WwlnWPNsZ
tq3LcPIaxlCzcOePtovrwPH5x6BCTZQIT0yeS/uVkLMKPMUt+kDfAq5gpf+wCz83w/ctI+oCPEZg
YKT0U+lmgmGE654uxc4//yXp4IZNnLByh8F42q3c2XYXnZt9fS891bDCg2KoqFE1FYtRbaqesByA
QcZOWWlUr5pj9SUGi92iKk4ksIVnvh+sSiR7kDofOMvP7YXRvzWHDShX6B1VKzEY3XgGUDJH+VNH
3c+14JwPzEQnZ1HdrtK/BzGsbe4XVMDttUjn/Kp88bL2UHymxkGapL/U1EilUIdtz3cBP3GsWTZL
kWq1/VLwfvkHnCUdkXKrW5R8hvrFdJ+IHiHeinfjw7mETaUQVgbQh7kJDil6bN7oZJm/br02v0/5
CiKWxTpQwJ9vomXny5NzkTlameCFWbGmF0hXAC/n2MVAYa4qFqW6KxowhcdPuQe6Jd0psyFTV7Ut
0m1aQSwzi1tNkY9XH0+Qn7itdfbAzx7whXSRJJJN5ZIam8V0ThqmPws1S1LcasfJkmTGew6jr1dJ
e4AVdvPN4QEebwRGAzRk0wAY1bEXpRpkRLdRTSc3UqysGaGfYkR1C/CVUy31qyKRX8Qn+0fgmpvq
PXC486hP00EEB1ni0ERvnWhXwYYA+eyzBbNPeO+FMJK5N4VPMKlhjZvtZ2SwSlMTwHtnaT3gZOkp
phrsI7ZyO1xeUw+BQ53GB8M3F6fo6iv8cG+3u105nimoR0mIZ4k+bs2/AAhNz4fITmzhbDf4Ao7l
uMfTf9BepnJKvI8BOVKcFXGE/dh13YguS7wqA7t4PORzyv4F9M3CLrgV1aZhH6xmqSILq63oOb4s
4SbJ5qAwnLwfSMQ/Hgh/JDFCbP7o1Ov6ScNH1qswsSsn+wmpsAuvQgo1GyVLTds+DI4uS6PlXlvf
7O5m4HmgSs9ypvhFqlOHvrY2i6x0x42pBKen3s9P0p28A/CdD6qRvgrzzNx/Y8YMna/rN3ZR6Tn0
PIVQlwmU0YMC7gaIPN6SYrjLn/ldtL0oMnqVqB1SB0lGmdq5OtYaLXGhgj79W1vCvfk4GwAv48m2
byzgDVuULKIZHFhQutE++Xs1XbFQ3FEsISlSRnRai3VAyJKHXf1gggG/rlIMBEWY/bCZSYJ7Ryqf
LjRSUCSiD+fVrlKD2ZhvolBV/eUa1lYe7Kxqi4iMaeLnf1x6Crgd9nBQmsjbLtewMHsdv7dC1ktR
+eme2BazXrJfy8Hm1bVk1Sekl+bMH0hWeNkh/de6DcPn4pkQfsVkwLm2JWSRn0N6X9WWazgDj8gf
aYR9Y6PFX82SIN6i0bwXX+vyWQAp3IOaDfWj9nZK+TXxlZq82G2FNF3381Alz1ePMgR47982fpjk
FjST8ha5aFEOhlM1MmLc9fA01scWQY+sSIH1yEePTylLsKR6GIHmwPTRvCEZqOjwIYTS7xDr5BMH
TI+rfclmtQvgJC0fFStMa5hDFVdmKgRMSFlU9877S8c68NpLG/ZiRTojG3DBfUqKX5Yw7YiP+Kky
MJAi1ODkhd582hz9JIybc4CAb0RbCuWbrDwiWw3NvYFlbndrPiB3+OA+HZScHhE4+ArvvNVObFFJ
Q4uM9E/gILQ2cSmMihwgtUYE7mSeEiBDbPPCLl+JUYnUBbQGwn1oxINiO8TuRDBEVv2861KxQayJ
vVIFV4vIbToL1u+jOIRDNXCQV+LJ1UkZXUekE90IOA6mab8+TT0jFEju0Ufo6T0340nGN5tAK+k/
xIspZktB1wVItrJLhKMpNEMcM7oqqJ/zq4kXKxiiwnt+tb5t8TcdC2elQBREJjY2i4TmSku84HC4
Zpasq+zoIbdh4U2WwYFHdptgxOs12mIk/fXbiXJMdhjttecRG7C9U1cj/eP93wvFl2jJ2HfWcpd3
nmAcXa6ymU64I96BzbT4o9z6WlCfIihN+kfnS5CkwCRgoa9QTxINNQLy5DN+K6D9TZ6OILTJ6CS5
x/Wdb5PPH8B2G1QoadPw7lW/o2LQSfhxpj8zrvXHnG86xPsBByuO9jpxJKIynDbbPDupSgOznaZq
QySAzTsHSFjtutBIz3MuL+nTIc23ykq/ANPuyVUPwfU7k6fkqp8+3ijBLsGK2OLjB4jrvhTMcuHn
Hmpq3uLIfAImTGvej2okM/UpmMbUPv9ncnaMkNEjlyj1gc21tabD0GAYeYCWOXP/861vlnMpVd0H
fWO9tQDzQ1/rEt/Cmkm+5UZZtxrGRdPbNOPW4BgrWEut4OAllnyzsG0i1DwVy5xE+jUwdciB2OIa
u7BzeVEGsacp8PeoytCuPpm/tQsa0UjVeXGB9UjmU+IzhuuCI/y1HywYDF2sXaZ5d/VoRkY+q8UI
dEkoG+QvHqcFX6mn2w+dROihOGRtlqurMwhwRDofypZ5kbfpFUikwmwZmF/J5OihKNer7g2qWRdf
1IIHG5EmSFwuvykjS03AoERwW1c8+MviLj0wsEnRWlo4adVsHDCIi8oxNVUSRUHCTUf5D4cpOtjh
QlkUqLd3UseKaAsEy7goic7fACIJzJMzStFIgTlJU6C0ARGqLVjAN4Ht56NrqwNQSlkiK29xy258
xmtPHZ/2vcTnUf8vEnhIPbiobt5crquAhAkDQ6dMZ8GKiVWpu9bhPI2ijeFxW1/OJIT9PiqK0EC9
ZGWFJNTRQO6s8xYAKPD7IYRBXzyvGZSuEHWGt9sVbL4/9lhs7cy8/lLwrh1FPsTtcbqiLudZj9KG
glCgxuk3KqtDeiCb7SG/4mL4/Mg01HOrq937ZmmBMHX1+VZQB9OXTl6fEOHQGXnM6iJBPDyfhE+i
0hzKnxr5ZuSquAvfJ2hoRI580euRorj+DjhSp5zakpDeC4jRyV/1ILm72pV0wFFOuHlKCPCVndax
vkcIlWbCY4Kxt//iYAp4h+HvIiyQmCWkVhDgUcU+t82X5rvivRlTDv7kwAqTzq706QJVkNN8LXLv
4onyQhl+lUv/ZAwnl0b4vGz8HQyuhcS7FdfWUvHdrJfgW7eNBlBiDMzpu4q7Heln+kx09ukcvYYm
bCfaTgGjBEVctP5fCYwPWJwcOnQ1EAtL+D+z5x9yV2f9d/LVn6/uVYB3QGSaROAeeExRbX3L8YMM
mxjzJ1FcbfAEb6y5TejqarEvDPcYxMyEldPIPIoLsWH9nLNdaIOBijZawc/yp3/JjfmYexFCuJ3+
FYfqgGF3G9DzD/caB62RnlvFU5wIMm/vhuq3cU3fflqITxFZpQ74zuvdOJZ2Cidw4tIL4KiGIryk
5YE+cZ8muNzOirX2o2+NZlwlLdR+3vj5Z1pX8N9wNHNOADjKRgU0cQafNDvmbDRXPHkiVLE4Sxax
xRXeydGDAfXlBXKGWBB8kEug4WR5xHkkNHvTPc7wWyO5wLlXSgSyUzd3hSrnnURZZVCDmnzwotA7
/bu2rORWF4VhmV4KReYzJ3juLOxJ7/B2Ggn+SvPdX7krTx9JM0aKabmPEs1shgGgkqDe93pAsTis
nMG/K3hLMztZtCkRQDKhUks9HTPD0E9G8EbD6X2JaXco8LV195fPQkvLZwxFY/Mv/ecr59qY69es
3TGSml3Q/Tz+UVTfwTRSncJnVIYnYA+M5H3Rzpl0RKCF6ggLulM5ein5obSifT8U52Ah8fbJgpH+
47I8iDLDrVeJb6+KKsEDZDxvQxpETh5BcEAoH4m7Ah6UYJ1ze/hBf0wArAZk2hEqi9bxtonn2gP6
BuhZ/h74BKRAw5621zVUxbg3MeLiEgYg+YyvbKYJQ/2RdOmVvmn0KQ2uzl/RClfTR9/gI+mX9cV+
SfTp7WE1Etil0O5a3/q0S4h5i0McW++R7eFnSWDyR61tLTanMswoZXX1IUQG4YsE10o3HuWjLU+P
9RVuEnCmRXA0/UA0wLAp63J0Y+/Vc6TOdvnVlMApQASEs50dGw5Q0MdTi8jL5OpT29D2/WcWokR3
lP2Ca1v+OcL7J3UySkVepXGd/Vp2oaTDe0CYWiNOoxDCxuYyu1DS0g5vqqI0Ti8AKF8gJnzIN6NK
peW1jtmqEHl2Bn7klMX358j1OMquYk2ccS/y8VFvcBMEpXX0MJ1I2m/fhU+GRYwMENn+jew2uVHY
qNK2Pl2LTdOZlCQpuXxUViUSny8C1On81tPuyRS3Bedx5YXlypNS8lDgIVNNIOTpusr3cMlPYiIS
k6LdgMKx/lTdraZwYiDM35Waka5uTDlfeCxKMJNLMZ5qPbTNFYYpHHNlJS9ToDTZak5y6XTUsRA8
4U0tI09kR9sXaJEON990RZKciCSOHZqB5Y/GToFUAdTqZ98YykaP5ODPj4LUjSS0fPwihsB6/ALw
Uc5De5VWmUeBDDvK4ucPpuZwzAFJyRP2ci1vRxFhmm1OKOrVV5I+1HpV4yyNRRQpxkgJk+c9aceN
z/W3R51YVSLMtOeqdT4DkSVX2TD0TG84W4vnLS8XRV8dONMO6E/rGTp2HaKe/qQAMfZN75dCsQXx
hK+R7mdRUBt6khNlf1F8MFZIx1WLS1O8PjFrXJghKQWXbtlHikelIuJb0OJTgzyQqNH80hVGc87H
sbqEYgWQa5gH/PstVlLJM7zqrExtgCB5Q6NGYIW8xEJOXeUGk595WIiMTdZTKSS4CSkn5z8zMvK3
bW18iK6w8p5gk+NhDEsHzRhkZr3j91liF0JMXs1IvPwFDKl3VSpW2JkHc+/eLRQ1/xjMkSldaiRx
Jkv0Zq4rwy2+izTCAKBflTlFoI48OMsxxtM+IduYzJdU65WhFHkcYsCdhzr8EZwMIoFNRhDA/RjB
TybV0P+m839SlpMWbspIWEOMn9CehNQVu/yIhrNI7b6GiQF1ZM2+Tb089hRC2uyOA085b81qd036
68OcnT3AFO+6cTCe89snm/CJJlPbYTBjhdtJF4U5qcpm024yv3xfibXbzKORL5/h555a6UAXDDc9
ovB2FcfglXL/3zc/ELUBiXvbun01tvrw15ZIzqu/6eDcse2fjz7kfeZ2ySxb5+8tTa90Ik40OwBQ
RUnkaHCGP+s3nFv3p6mDNM8tYsH8Y/hFJwAVJ51gIH3YUNnBXUc9UkdhFgd88bVBtsbv2EKHnsje
Kpigesm3SJIe4zu5SoUU7G1SQFEsaSvRsrEz77MExGGqvtPu1Jl5eC/CHZgfX22s5jgGGjWTtUIh
pweAwQKGhbXnC8C1LveqwN3I/IXOcJX3cqTyaQwU7IsvvNU+19bZHBFKhCj5louZUDYs/GUZ1n4+
iH8seZX1scZwlOqS2NXSHQkBYMD1aOlNY5UHzoiGYwqSuUw8/om3xhr+fMHy7fGASVk3CSWEAyc4
uIOn+CUVUTeo2L6vd+RJuQoj0+yzVyh1gyxBOyT/gkbkN5WA9slF7wVfGljvbGV3LdhLTkAx11hU
zSi+VRuW0acKW/xH84BSAClbV565YQuClcfrPjOAg3GEzKiZDx2NZfhup3k2msc9WTSKm1fBm10j
FLbsxCihluxALtn87rx6tahbIUj+hl8p+dnm5nhrwjdQystC13KOhTzdA0NCimA0C79ZgvtyYa6w
j9+Uqqx/1hPNXqo3wcCi7HcaDe9TNOk6KjsZyqX2DRrIf9bvblrqGDADNkTIFlDEOYxPBqG6RiBh
MhwILE3UGtm0M90ZQ3UnBjjqX8d2IXRnIryJc3WGXf3o7axb+jk2PJALn1T9qw/+An/09l+ychGZ
PjDsawxEtlBjbu9GbE9RDhaY1PpBHpM8reVtZpVcSkyBJ1eI9D3ncfQW+V3u1cZPNOhFss+iBM15
5CtbD88j31SZ9UbcQ8SyPd0Xg7YtuaMnor99ndUAe8mfbRUVL6nQjq/89YaqbPntFU/klaueR71m
6LocSAha6SBBKstiKab34hxgtgZrb6YA1a1xg8P17rPtUhmqZSp3UHYdbVF0836botbDRZZYlIrN
Sb5DKHWUF+OgrALfafTGj/YmmsC7GjmEbNHNwjj6bSnhk7pcpBVJxsF63y6A+L6v8jbDkvN30F51
WH9mEWtrjzSoCy0CVU08jwA1O58Y4liePEbIsewSOQRsmdSrZsUl+a1Kv+PmAggXSvNzujw/4T3b
BuXzJTFpzGT3eBSCwuyCOtVj4bFg2e7xbf7A3f6+z5ThtlPIO2yUorCyx4/0fEgoyPJRq1ABWGCn
aUS7nRWyM1j2q+OB5fgorkq2ZOfu1HrTH7etvC9UK2slj6eE3GWiXOpWpyN66ZtgCLLhQoq4Zq9w
mh2meRGGjaIvtYpL8duCxLYFO/CG1t9sTYvIes4LLpJRLMHnPqyNdYRTCeypTlgtZW65AGpwUbUr
Z7kNoZvUzPBsSTu9qZUUi1MDkuzq+UVvErKldM27GP8GBEnBZKtdmxFOGHG5xsJnMyCxFLEb/GFV
RYo6Us7P+cX25m6fsYFL9rtTSAbFZ5csdR4q8mdxuSxT+gCwJbmVtEB+k9JnIIksQOWW73KFt5Zd
IdareKAJhKQ6tYeBNptIAONRyEJRGJlDUJWDLPUUTeofrwICJPrLiWfj+TOWh8TeodcUYkcjX6Dn
Ie3t5yGIphbTvq80+D6GIPyDRnjAmzBBIN5Noe7zeDTBHo4hd21iUwKcde6X/xnMtJ53gbZWny+m
3xNxfGlyXKp69GWymTP5iluUww6MpATyKNaOW5zw310w/yqkmQuslLczSy7t5kgfcDTeDdqkpKY/
RnvIB8YNkhrZiSQrYWxzR6uQ1KKEmDqy7Tj03m6zjfnT48Z7FsBKhdwwlt07v5BuESDu37a50c/w
bilM90rHmM296TiFKskZo9Lw2qENH5E+lipGflBlZ2Yc6Z5/tFkRCiIMkXLl3pE6kri82na7XRva
rqvYLjSmFv/gxuFHa9ZwTzTlzgAVyTV6Tri/74OD3Orl4ENxT0RBOf243ugEdfwUHTK1SkHZkan0
QU7wKMl3nZ5NGzeY1ynd3F2fEeLkiA5ODyiDHVmBQyycoYTCoBE8OlKnhJArxdcqEDECmmVVZxgA
Lb5N+qcXNOIL39XZaRSWAoRoVSUkRp9RWi+U6CDy1iETZ1rvwHxCUoM0eXtkdox0/3lLwx5pG4OC
Bpk4NsTDpfjdBcFvcXs1lFsMkKLuGR8qi0OTI6vR4T9S61I9MDCXD6e8zgkffO+Ls77dK/1p1gjk
kFzmQmLa5Q/YO1P5Q9s5ExZw0Bb478MpKYOI1BslJdhWzmHTfr65YhUAZ8RgNFyOFE6wavsvA8Nq
Q9n2o8DY1b1FGd0oLkqp5pavjFFtJhXeiGoFGfsqRCqS55Z3CLIqqb1F/SP/ZL8rY6Q8zNdSzllx
Qkd/sGu81n9MoWhETCrsPI9uSrSX57bRpQT0y+L5SWWHkAOVoixwju6wMq8CJzwMazl9crFC4WCG
VfW1NGNbb9QC3YYDgfVT/X2q67AKmgetIOmZjvAsMy7enLmQui8oMCQQHF3ri+QdWN55MyO91Dl2
PeHR09ZeTSDXVLcDamiGoZojfE2foUbeLehnbP/DEJ8HFi8WxVzNsjxZzWsQaMOlxzrORoZi/nkV
rWLRFh28+LmiFWn5oWD5WcpFlOQS7GsN+EGi/IWiPEOrU8WO8ccdvBE0Ee+iBZ/mT1j9ewLWU9XC
6h1VnqTOlSrHI8fqBCHkym4jS+UYWgVow+fdVjGLKzOYJMgl2Gul7rXmWq3T7/JrA/mlCCHOsDN7
xNW28JfqijD3bk02/7hmInJJLD5QXPAeIAZHO3OJ513uJpgQAIsxmsRgTrQwI5aOIC8ZyYLWyoub
j+a7Hju3UgUGcrmwyQCp5sDxNPnK7+n1VyPysKgcjSZjazU+X0LVr1ycSyCDm141+C4yJTB+vK/x
qHz/Mr+WTC1SJobd6KRscKBqnNXa3FhJq8SgtsnIsdlPlUlAsuq1/RZNT0e1IcwN6/U/b+QenSc6
ps45SQc88QpduoLPMblCuELUQjR8Q2PGBbqzNBL83PhSmksp2Jux0PHvHliHKebl+T/0B0q+CEQG
nO5f71Fi2yNvML36SC0bA9UZu3bhFjY0jLD19LDpH7rlbh/n1DuDy7qM1Ay7RkzgwL5aIyUjZHaC
yOnwe2dvJ/QvpxWt67JIRv7Vyf8r+fWSOzzwQDP2MpxO1g8yGbjkLd78sQ+7guHWvMhtC8a06Ml9
EbPoXTsdZ136T7lRetMCrGIox5FjjHY823rSuWajpku3HGBSqRnj8YtSBJXF6FY5ttly9ttsm3TT
LSl6cVLDxVWo6sxKDd/Dblb0soOtf4uS9tnElUGaSHLhrBNzym6j02ULSyZJ5gehitUesSVcch+r
tPBVuO/BHwKkd+46nwZrj+W2IXY1lnA4LjD+WpfYJrSTuZzhM3Kk2oyeJkqVlexQvaOPBzalYS1b
MdvyvKHpYJnspn2cScGWESEoq7s7YBNwt6sfwjyFrxFCPq9AMJuFGd+WgVtLRZwQwCBXz4H424I/
ppPHJRh8bb7kqVhiP5GNVpUGhRo+Md7FWigzgFAhXh5NXPHWzOMZNh4kGenhxmbLUQr93MEbl4C5
QbHddqf1MF0DN8IRJbNE8ZFUPpWjhLw0+EeDa19a5WJeKPyvb9MylEI7eXpbZd5xRUqqNyq1zFLO
VhjcauRbRy4YiuzEsuoa+FzhN2rZ6rnm8Nh/4mNTYvrD/UyJCaYDB0M+7fk8WNxYxBr/2wxteVP3
S3RnMAUTMLlg3dEGVcxNZs0nehRq/hAzp2kSpJrcExO6HlQfWpZOcleiXWUHcVow+uKxEUvvmtsl
W24mD52qxz+BFeBhjt6bKHxnj8qolmcfrepjuIdGJyve31s3PgQSCAIpMwUF2N0mzMI4QuO49+jA
1Obkx0Z2XTfoikB8jBdINeeQocJ2PrE0wPjoeOnk95IGGR2kjf26++EeMm663cOiuYXl/On/UjHi
yz/hqdZsdZ4TWjlYDVnEJwt0r2diN3EydCbUBjT8pTt9IpoXgIDn+Kqn2utyRVHLTZs2nACqKbEV
Q9/ADjIxmla6A5fgzAQeVn6y0EL3KpZf/8xt5zkAN1HCNabHzbLp55B0/7hKCDGlI9yrdQ8C7jDn
TGj2JcsN1Nvr5RDCubP7S5JEoHg+PXV6HedB5zQjG4eSQGTCN+PnMQH6yGADnVFU1z5caZCaNvsM
FJ8OcZV0stpAN9ChURdrusnbWMWY/2PWL51mBLuKP7+wPITuYzA/oVc2lc5QwS8fOVkaB+73ukIK
keX/eNcL4NIHmZmiTmirB0qzUI4min76RXrr4eMuIFCZWgDnGcQ7oUDsda3OGZWierrzMATl0OnA
jBVJ1cg+DM0D9E3/maz1VH/hmAUeWEQgX1pOVilrC0wniXVZ7CuqqkIPx8ZhRcY00oetCObNxEkr
E+pATEsxvN2mhjjZCc3C2I57sxx8C8mjetOYaqUWOvFEe8eaq3bGyhN9bOkt37qkXXVrFOS7rGdf
dD3ESHylygRrZQjRN64g6EAEolF2mxnqVhRWbhGnQWoIeKlVjhWFERbhOZtn9v41u3D4ox0dlp3t
raPK5lKfsTD02Lbq8nKF6/SZ5YbcLUOylYJxKnB1MN/9di2sMae3Y15wms8oRKkzPlbH3fbuzpWs
RkYABEJ/MV+Oxzpk/ega9UFnoXGedg2P5mctmet6egh/duMGQ1ZLmijuLPRL4fN2ocsXgNzVYLDx
ovPPNkeVQi3277mRUnsD5ihegmWGcp6UGJe8ijUaT35V6IwZ7sBneqtUDlAlzKdtNbPyUYCKA4bS
ruDuImuwnejczzHQ/Hin4/J8NYiYx+V7zYR9+aBhB3nEuUabK72J2vu5cE/F4dmhtlCnHOdS1hUX
bFiFnE2ZBJXuHC+axatqkTyPytYB6qe12kpyZ/MC31O9Ky0sOmIFBkFvRT2+ZvSmeGI1a4ppo/kE
7nrwQ00bzz2PH1Z7ZTvU2RZnavw/nqKDLGLGcouUvB/JvwdIDnSU/NM6wDcNc9jGGbH+erHz3BTm
HCPBBAaaDbVuiJRxREYp4F7/WpMD6PQs9NOHdSuVSIg8+/gjs4g187Oi009iNpUWEy1xuI64rjRr
ZkXdlpv+yRTUdjjqNztHo/9fNHEtQqGIp5AwR0q0uAJm0gAeeNiofAfpxts9fYbqL5jwqtS4D6Xn
onMIabgd7GXxngUSVAgib7dTWDiOOQnjWAw7X6LsJSeVPzORtl8SwBeHxsmo0FtummDTHeQepvaN
+2ruhtKRdLhRNwBDUG75DOgIby+4KJCTK3oBqsVGdXTiOL7hFgdE1KTWhWu2u7WDzVYZbktzmKeH
kkrQh6lr6T2F30TWnQKg3xI069j3x7X/tgvdvoIxdEu3Yp2CVGC312iK/xQ8hg6cPu/EZMrQJO19
S+s9COTOmSjo1pSWt85YHYdVBc6Z2HXBh0+wSIN7wS6PLttV0rNdK+l8aD5zeiUWhiO4lhJAFe2o
OcN26dYDEDQMj+ZUacWKuW9XKftoyWZZyYN2r5cyt2TIsETIyjITqYdDvrV+NkYKlt1bCWvdViJ4
5TLbzSSuzLtUcu3bBw/FpG+cHRxM4V5yyELQ+65D8qtzKc7hdLLbvKxxSJRdgyNneY5uDUFPj8Q1
cA3G9Gxqd9ND73tNE/9DHM6KqcHnFXeE2eMB5Mx2u0dr7aMJCzn6Pt1EtzoWuaUQzZyzKXAXLVXz
Mvxs6KIiGGvYQ6lEQSazLYTKBrWEeFccYNzv8Sa8LLRYXNlKVq4LtNNmpebsejOMKpHG5ZTmeubs
SkfakFZXwHIJo99Hiz1VLnkd4TrY0MXHGSFXcz9Ncv3VjjI1THrPPOsudsZugmucHCGAx1VROFTw
H7LVzjE89gFRqo4ns3PkzGg1NXrDmP2mLQ43TYu310uPtrBFLKAs0mJQiC0jaAkhg9a0q/OGsDyg
VdbE8mX+GvdY1bnJOZqyu0M//5Lq4YawevdXDmAcVo22LJr5I4Lg9Af5cPE3BI5VXTQlEI7Ik7HD
2G+HIgs/vUOouytaSYfQ1U19OyJlcGn3nHao8i/bBD6iDaOOuna5hZwbuGdkVcu7bfvtcEuXWyyP
GWp4T0H9LP645D4JJP8CQaR5RBi43ZY622dCwr99c6RE0Vz7SzcZYTQacfphUB2Qwyj/ike2Fzxx
Nnw585muD6s45iWlLVAsTlglNyhnWBRFmfbIo2t7Zb01C1neO9lmsqBiN3xwNt/EiwRtYZX84G0l
YbBqxhn3M+yZcEjt3l7GS17tTWfkNGREuTV0ae3iCsvZARv0886Gxcv1+f4gCvSNaSuVi2rwHy1r
ZUDqnGSGo51inc4yAbbq5zCAsPgu2lr9NcAXvz7RSSFzRiSMmjb16GVAPs7NKb6ElOEfy/et8egM
UoveS8h+kbGPMXUA97NylTJpytnGnrMR43RSpKL6Tq9KQEmUJnUbWO1N/yI1wpeg/6OG47f5l8AF
3/2JSJdUJXA0CJDBMQRHixHQLlx4I4/PFhsAMeZZgbhxTHqUiU+pswP/7GGoO7vG/0v1pcZBpfB6
kF/oLljk7lf18Mg9UpIBzvBkNMXhb0nhpD8FqaO9DxTD++BI1D32pD9cBOrqptywxgk7UkrK6zID
qEEO8f5LHD4s5ygDe8WVa7BmLHaYooy6sPbIPpOesROqx1TuAKB+jU96ZIz+/djX82lLrQzuXtHt
2mPNNJwqYLdBiGVwM14z8A+Ul3lRi4GAo1wzI31WRFk9gIYQQZEGAhWkpm0WKH5N1rqJJToJm//P
i5HSrTTkjqVgjL7wU1eDD5N5ppneKDRExPmcjuLrln/NGOO9slMqPhEzB+oqkXQgRRBl3eTCUxxB
4vJfpk6dyi033aUrv7uK8ak5XrC31iDXtXRiwOyidGh/NaOoXMieIqc+c3mBVrR9G1ZKZ7Tr84rD
7Vh6x2PpsQn/gFLid+E9s929UxK93ZMhljn1Sm0FqAfY3oTz/Spqy4UE9dw78ZR2+xxCPke8Gk1J
XyjdFnrLClKUgAHTw6iBCzFytk0oCDoCGzhNu1pnPinELbR3QN2EUIEwmim6+TfrDttc6wLW2lL2
/4c+q3jmcE619porIpW4VgF11fZKU5F/CjulsGx0X4cs0jNKgNTYp0nxfTvD6XcTnXhkUv8Dt6Xt
2Yya57T6CuHA6rfrT7Y7Ns56C3MjOAslkCpnyM89T05aSbPiMx6GjlgIyba74NQ0tbccHZqxbZoj
4gR01Exx19qNdA3JA9Zn8ATI4yjNrqq+BLDfBJ0yvgFOosSwAyshK8CNey39+h71+OSmxcl7dvgp
33+7CyXrK6rEBZsPK/gp1UYJPLsm78o5T90jalx8bXVLlsfjD7H8NDkITmh4GYlw3D3+3lzmharC
7W5tVHqUFd5vZCjxGBhE15IG1KvJNStfeqSLy3qHvIvMhAvlw4OL3CcVgxu0EkL68c/M7GVOPwWk
tsSNpvd0ZV94df5/g5OrrDV+k6txnbFOOICNfYda0swtUFz1j+MCtfvcvQAFbXsYGbIgthd82KfA
sfwzLKKI7fh6GuNGTmfvxOH5rIpgpz2xiUkHGm0fk4M2VnkjC/gLah4ezK4PeLvQua3x0qvcm8u4
iqo2tziz+N4gVZcVSsuI4/QSRGVRqWUU+6ywND0njJfG0FVERDwkWR9lrxDv2h+m0mVqKoJG9uRL
1d9QTt2B4WDHLxGF+YDXjuI+/8w2TJhOaKmqiynVqCrXoUCSRpbOkVGvN6CzUZCJkha9ycjgNFNe
ofNnxy3knTWT3PKjNw7iJ+9Dy6ZeCnEqqiDrsxLQdEQSpIag4OMBpz6NwUm4DYwv3X3hbhzZvFDH
bBikUj0NfJ+HYZxTeN+IU3UwG/rIZIqHAeXB60b6XxBJdy0CllBK4dVkQVgSdLriyfNiSDRq1noT
J82gta80KHJkN+/GVN3Bo9OpEb1Td7y5q8C9sNV506WNb4Vj2IJN1mn1IchNDrLCfMC3n/Q1/gjS
oEn1RBZIwVcgwoPxIT7UgvUWdnBXsHVZLIx9ZnuYa8lmTyXo9kb7mOiRmkqwmd4lnZ9pqMRN3v3a
OFzmE7/EMa7Ns0GoTOK0t8YnfZaEiFpP7WjXfUe375jgxQEekuLdtjS9crl9Bj1yvZGAl1VgC3lq
tummiuHXs0T9HiOwRPad5a4DB51HgudeaIgr1kyFiXKEN3oVmD8tC8jABgDqlcqaSkymxFURHg8h
T4+/+2LuhjpKCCNi30E19zR0kW4ju1l38U4hM5yJquO8K5q7nM83KYZu0YDJUerLOq56gUpnmUZY
daD7+kb6x26b9aEd4cFXBUNRHaHZ6hBxVt8yDyD0wn2yQLJb1NAFEcGxjuPqOFpZ87yxSNtlQCyZ
9NOlbFPrl03GG2RiiAU9x2I38tPibgXh4KvSpSQK1ue1jqJEj0IfHQcJHC7iGEad4HCe7+bmcQWt
l0F2U9lS0TaILY3p6vewc2DnFNHFrQULk0wEvtFJ48VAwz/iKSTyrtIQgaqzlrqz6Dl7hub/1oM/
/1gNZOJ1ak1jKbu2sf+xEl6obYysJebjFbL+TMzFzhAH44wm/CzbL7B0VVjoa0c6P0HjqCiXaEtY
dydrdvYj/YWxp6DrUbqmOjflD4wvh7xp3NiRrqFGk4f/HqMloKHPbWf19SLvem9H0ja/FBbK8Tag
yECFzVaJObxCM8MJQ0NARBA/dr9xQuMRf5FQJKKzAybHe1A2It5R4nl+DRv/pHC+H8BuuzNbXzSV
wUojI+/Q61JbMmcJstPMaUHZYY/0wbBgDLYWs/z/6vOeVlVjg4UzB3BXXFAOdnVxUZJyca7OedF4
REVabpqNnWBY6U+qUO/1Xnmo9VMKWZcO95eFnbsYaZKc/J22vlxcV5W8PALqo8D+WkpJwlyFj5OZ
NMvPZEkJlAU=
`protect end_protected
